// Copyright (C) 1991-2016 Altera Corporation. All rights reserved.
//  Your use of Altera Corporation's design tools, logic functions
//  and other software and tools, and its AMPP partner logic
//  functions, and any output files from any of the foregoing
//  (including device programming or simulation files), and any
//  associated documentation or information are expressly subject
//  to the terms and conditions of the Altera Program License
//  Subscription Agreement, the Altera Quartus Prime License Agreement,
//  the Altera MegaCore Function License Agreement, or other
//  applicable license agreement, including, without limitation,
//  that your use is for the sole purpose of programming logic
//  devices manufactured by Altera and sold by Altera or its
//  authorized distributors.  Please refer to the applicable
//  agreement for further details.

// Generated using ACDS version 16.0 211

module max10adc (
        input  wire        clk_clk,                              //                      clk.clk
        output wire        clock_bridge_sys_out_clk_clk,         // clock_bridge_sys_out_clk.clk
        input  wire        modular_adc_0_command_valid,          //    modular_adc_0_command.valid
        input  wire [4:0]  modular_adc_0_command_channel,        //                         .channel
        input  wire        modular_adc_0_command_startofpacket,  //                         .startofpacket
        input  wire        modular_adc_0_command_endofpacket,    //                         .endofpacket
        output wire        modular_adc_0_command_ready,          //                         .ready
        output wire        modular_adc_0_response_valid,         //   modular_adc_0_response.valid
        output wire [4:0]  modular_adc_0_response_channel,       //                         .channel
        output wire [11:0] modular_adc_0_response_data,          //                         .data
        output wire        modular_adc_0_response_startofpacket, //                         .startofpacket
        output wire        modular_adc_0_response_endofpacket,   //                         .endofpacket
        input  wire        reset_reset_n                         //                    reset.reset_n
    );

    wire    altpll_0_c1_clk;                    // altpll_0:c1 -> modular_adc_0:adc_pll_clock_clk
    wire    altpll_0_locked_conduit_export;     // altpll_0:locked -> modular_adc_0:adc_pll_locked_export
    wire    reset_controller_0_reset_out_reset; // reset_controller_0:reset_out -> altpll_0:reset
    wire    reset_controller_1_reset_out_reset; // reset_controller_1:reset_out -> modular_adc_0:reset_sink_reset_n

    adc_altpll_0 altpll_0 (
                     .clk                (clk_clk),                            //       inclk_interface.clk
                     .reset              (reset_controller_0_reset_out_reset), // inclk_interface_reset.reset
                     .read               (),                                   //             pll_slave.read
                     .write              (),                                   //                      .write
                     .address            (),                                   //                      .address
                     .readdata           (),                                   //                      .readdata
                     .writedata          (),                                   //                      .writedata
                     .c0                 (clock_bridge_sys_out_clk_clk),       //                    c0.clk
                     .c1                 (altpll_0_c1_clk),                    //                    c1.clk
                     .areset             (),                                   //        areset_conduit.export
                     .locked             (altpll_0_locked_conduit_export),     //        locked_conduit.export
                     .phasedone          (),                                   //           (terminated)
                     .phasecounterselect (3'b000),                             //           (terminated)
                     .phaseupdown        (1'b0),                               //           (terminated)
                     .phasestep          (1'b0),                               //           (terminated)
                     .scanclk            (1'b0)                                //           (terminated)
                 );

    adc_modular_adc_0 #(
                          .is_this_first_or_second_adc (1)
                      ) modular_adc_0 (
                          .clock_clk              (clock_bridge_sys_out_clk_clk),         //          clock.clk
                          .reset_sink_reset_n     (~reset_controller_1_reset_out_reset),  //     reset_sink.reset_n
                          .adc_pll_clock_clk      (altpll_0_c1_clk),                      //  adc_pll_clock.clk
                          .adc_pll_locked_export  (altpll_0_locked_conduit_export),       // adc_pll_locked.export
                          .command_valid          (modular_adc_0_command_valid),          //        command.valid
                          .command_channel        (modular_adc_0_command_channel),        //               .channel
                          .command_startofpacket  (modular_adc_0_command_startofpacket),  //               .startofpacket
                          .command_endofpacket    (modular_adc_0_command_endofpacket),    //               .endofpacket
                          .command_ready          (modular_adc_0_command_ready),          //               .ready
                          .response_valid         (modular_adc_0_response_valid),         //       response.valid
                          .response_channel       (modular_adc_0_response_channel),       //               .channel
                          .response_data          (modular_adc_0_response_data),          //               .data
                          .response_startofpacket (modular_adc_0_response_startofpacket), //               .startofpacket
                          .response_endofpacket   (modular_adc_0_response_endofpacket)    //               .endofpacket
                      );

    altera_reset_controller #(
                                .NUM_RESET_INPUTS          (1),
                                .OUTPUT_RESET_SYNC_EDGES   ("deassert"),
                                .SYNC_DEPTH                (2),
                                .RESET_REQUEST_PRESENT     (0),
                                .RESET_REQ_WAIT_TIME       (1),
                                .MIN_RST_ASSERTION_TIME    (3),
                                .RESET_REQ_EARLY_DSRT_TIME (1),
                                .USE_RESET_REQUEST_IN0     (0),
                                .USE_RESET_REQUEST_IN1     (0),
                                .USE_RESET_REQUEST_IN2     (0),
                                .USE_RESET_REQUEST_IN3     (0),
                                .USE_RESET_REQUEST_IN4     (0),
                                .USE_RESET_REQUEST_IN5     (0),
                                .USE_RESET_REQUEST_IN6     (0),
                                .USE_RESET_REQUEST_IN7     (0),
                                .USE_RESET_REQUEST_IN8     (0),
                                .USE_RESET_REQUEST_IN9     (0),
                                .USE_RESET_REQUEST_IN10    (0),
                                .USE_RESET_REQUEST_IN11    (0),
                                .USE_RESET_REQUEST_IN12    (0),
                                .USE_RESET_REQUEST_IN13    (0),
                                .USE_RESET_REQUEST_IN14    (0),
                                .USE_RESET_REQUEST_IN15    (0),
                                .ADAPT_RESET_REQUEST       (0)
                            ) reset_controller_0 (
                                .reset_in0      (~reset_reset_n),                     // reset_in0.reset
                                .clk            (clk_clk),                            //       clk.clk
                                .reset_out      (reset_controller_0_reset_out_reset), // reset_out.reset
                                .reset_req      (),                                   // (terminated)
                                .reset_req_in0  (1'b0),                               // (terminated)
                                .reset_in1      (1'b0),                               // (terminated)
                                .reset_req_in1  (1'b0),                               // (terminated)
                                .reset_in2      (1'b0),                               // (terminated)
                                .reset_req_in2  (1'b0),                               // (terminated)
                                .reset_in3      (1'b0),                               // (terminated)
                                .reset_req_in3  (1'b0),                               // (terminated)
                                .reset_in4      (1'b0),                               // (terminated)
                                .reset_req_in4  (1'b0),                               // (terminated)
                                .reset_in5      (1'b0),                               // (terminated)
                                .reset_req_in5  (1'b0),                               // (terminated)
                                .reset_in6      (1'b0),                               // (terminated)
                                .reset_req_in6  (1'b0),                               // (terminated)
                                .reset_in7      (1'b0),                               // (terminated)
                                .reset_req_in7  (1'b0),                               // (terminated)
                                .reset_in8      (1'b0),                               // (terminated)
                                .reset_req_in8  (1'b0),                               // (terminated)
                                .reset_in9      (1'b0),                               // (terminated)
                                .reset_req_in9  (1'b0),                               // (terminated)
                                .reset_in10     (1'b0),                               // (terminated)
                                .reset_req_in10 (1'b0),                               // (terminated)
                                .reset_in11     (1'b0),                               // (terminated)
                                .reset_req_in11 (1'b0),                               // (terminated)
                                .reset_in12     (1'b0),                               // (terminated)
                                .reset_req_in12 (1'b0),                               // (terminated)
                                .reset_in13     (1'b0),                               // (terminated)
                                .reset_req_in13 (1'b0),                               // (terminated)
                                .reset_in14     (1'b0),                               // (terminated)
                                .reset_req_in14 (1'b0),                               // (terminated)
                                .reset_in15     (1'b0),                               // (terminated)
                                .reset_req_in15 (1'b0)                                // (terminated)
                            );

    altera_reset_controller #(
                                .NUM_RESET_INPUTS          (1),
                                .OUTPUT_RESET_SYNC_EDGES   ("deassert"),
                                .SYNC_DEPTH                (2),
                                .RESET_REQUEST_PRESENT     (0),
                                .RESET_REQ_WAIT_TIME       (1),
                                .MIN_RST_ASSERTION_TIME    (3),
                                .RESET_REQ_EARLY_DSRT_TIME (1),
                                .USE_RESET_REQUEST_IN0     (0),
                                .USE_RESET_REQUEST_IN1     (0),
                                .USE_RESET_REQUEST_IN2     (0),
                                .USE_RESET_REQUEST_IN3     (0),
                                .USE_RESET_REQUEST_IN4     (0),
                                .USE_RESET_REQUEST_IN5     (0),
                                .USE_RESET_REQUEST_IN6     (0),
                                .USE_RESET_REQUEST_IN7     (0),
                                .USE_RESET_REQUEST_IN8     (0),
                                .USE_RESET_REQUEST_IN9     (0),
                                .USE_RESET_REQUEST_IN10    (0),
                                .USE_RESET_REQUEST_IN11    (0),
                                .USE_RESET_REQUEST_IN12    (0),
                                .USE_RESET_REQUEST_IN13    (0),
                                .USE_RESET_REQUEST_IN14    (0),
                                .USE_RESET_REQUEST_IN15    (0),
                                .ADAPT_RESET_REQUEST       (0)
                            ) reset_controller_1 (
                                .reset_in0      (~reset_reset_n),                     // reset_in0.reset
                                .clk            (clock_bridge_sys_out_clk_clk),       //       clk.clk
                                .reset_out      (reset_controller_1_reset_out_reset), // reset_out.reset
                                .reset_req      (),                                   // (terminated)
                                .reset_req_in0  (1'b0),                               // (terminated)
                                .reset_in1      (1'b0),                               // (terminated)
                                .reset_req_in1  (1'b0),                               // (terminated)
                                .reset_in2      (1'b0),                               // (terminated)
                                .reset_req_in2  (1'b0),                               // (terminated)
                                .reset_in3      (1'b0),                               // (terminated)
                                .reset_req_in3  (1'b0),                               // (terminated)
                                .reset_in4      (1'b0),                               // (terminated)
                                .reset_req_in4  (1'b0),                               // (terminated)
                                .reset_in5      (1'b0),                               // (terminated)
                                .reset_req_in5  (1'b0),                               // (terminated)
                                .reset_in6      (1'b0),                               // (terminated)
                                .reset_req_in6  (1'b0),                               // (terminated)
                                .reset_in7      (1'b0),                               // (terminated)
                                .reset_req_in7  (1'b0),                               // (terminated)
                                .reset_in8      (1'b0),                               // (terminated)
                                .reset_req_in8  (1'b0),                               // (terminated)
                                .reset_in9      (1'b0),                               // (terminated)
                                .reset_req_in9  (1'b0),                               // (terminated)
                                .reset_in10     (1'b0),                               // (terminated)
                                .reset_req_in10 (1'b0),                               // (terminated)
                                .reset_in11     (1'b0),                               // (terminated)
                                .reset_req_in11 (1'b0),                               // (terminated)
                                .reset_in12     (1'b0),                               // (terminated)
                                .reset_req_in12 (1'b0),                               // (terminated)
                                .reset_in13     (1'b0),                               // (terminated)
                                .reset_req_in13 (1'b0),                               // (terminated)
                                .reset_in14     (1'b0),                               // (terminated)
                                .reset_req_in14 (1'b0),                               // (terminated)
                                .reset_in15     (1'b0),                               // (terminated)
                                .reset_req_in15 (1'b0)                                // (terminated)
                            );

endmodule


(* ALTERA_ATTRIBUTE = {"AUTO_SHIFT_REGISTER_RECOGNITION=OFF"} *)
module  adc_altpll_0_dffpipe_l2c
    (
        clock,
        clrn,
        d,
        q) /* synthesis synthesis_clearbox=1 */;
    input   clock;
    input   clrn;
    input   [0:0]  d;
    output   [0:0]  q;
`ifndef ALTERA_RESERVED_QIS
    // synopsys translate_off
`endif
    tri0   clock;
    tri1   clrn;
`ifndef ALTERA_RESERVED_QIS
    // synopsys translate_on
`endif

    reg	[0:0]	dffe4a;
    reg	[0:0]	dffe5a;
    reg	[0:0]	dffe6a;
    wire ena;
    wire prn;
    wire sclr;

    // synopsys translate_off
    initial
        dffe4a = 0;
    // synopsys translate_on
    always @ ( posedge clock or  negedge prn or  negedge clrn)
        if (prn == 1'b0) dffe4a <= {1{1'b1}};
        else if (clrn == 1'b0) dffe4a <= 1'b0;
        else if  (ena == 1'b1)   dffe4a <= (d & (~ sclr));
    // synopsys translate_off
    initial
        dffe5a = 0;
    // synopsys translate_on
    always @ ( posedge clock or  negedge prn or  negedge clrn)
        if (prn == 1'b0) dffe5a <= {1{1'b1}};
        else if (clrn == 1'b0) dffe5a <= 1'b0;
        else if  (ena == 1'b1)   dffe5a <= (dffe4a & (~ sclr));
    // synopsys translate_off
    initial
        dffe6a = 0;
    // synopsys translate_on
    always @ ( posedge clock or  negedge prn or  negedge clrn)
        if (prn == 1'b0) dffe6a <= {1{1'b1}};
        else if (clrn == 1'b0) dffe6a <= 1'b0;
        else if  (ena == 1'b1)   dffe6a <= (dffe5a & (~ sclr));
    assign
        ena = 1'b1,
        prn = 1'b1,
        q = dffe6a,
        sclr = 1'b0;
endmodule //adc_altpll_0_dffpipe_l2c


module  adc_altpll_0_stdsync_sv6
    (
        clk,
        din,
        dout,
        reset_n) /* synthesis synthesis_clearbox=1 */;
    input   clk;
    input   din;
    output   dout;
    input   reset_n;

    wire  [0:0]   wire_dffpipe3_q;

    adc_altpll_0_dffpipe_l2c   dffpipe3
                               (
                                   .clock(clk),
                                   .clrn(reset_n),
                                   .d(din),
                                   .q(wire_dffpipe3_q));
    assign
        dout = wire_dffpipe3_q;
endmodule //adc_altpll_0_stdsync_sv6


(* ALTERA_ATTRIBUTE = {"SUPPRESS_DA_RULE_INTERNAL=C104;SUPPRESS_DA_RULE_INTERNAL=R101"} *)
module  adc_altpll_0_altpll_nc92
    (
        areset,
        clk,
        inclk,
        locked) /* synthesis synthesis_clearbox=1 */;
    input   areset;
    output   [4:0]  clk;
    input   [1:0]  inclk;
    output   locked;
`ifndef ALTERA_RESERVED_QIS
    // synopsys translate_off
`endif
    tri0   areset;
    tri0   [1:0]  inclk;
`ifndef ALTERA_RESERVED_QIS
    // synopsys translate_on
`endif

    reg	pll_lock_sync;
    wire  [4:0]   wire_pll7_clk;
    wire  wire_pll7_fbout;
    wire  wire_pll7_locked;

    // synopsys translate_off
    initial
        pll_lock_sync = 0;
    // synopsys translate_on
    always @ ( posedge wire_pll7_locked or  posedge areset)
        if (areset == 1'b1) pll_lock_sync <= 1'b0;
        else  pll_lock_sync <= 1'b1;
    fiftyfivenm_pll   pll7
                      (
                          .activeclock(),
                          .areset(areset),
                          .clk(wire_pll7_clk),
                          .clkbad(),
                          .fbin(wire_pll7_fbout),
                          .fbout(wire_pll7_fbout),
                          .inclk(inclk),
                          .locked(wire_pll7_locked),
                          .phasedone(),
                          .scandataout(),
                          .scandone(),
                          .vcooverrange(),
                          .vcounderrange()
	`ifndef FORMAL_VERIFICATION
                          // synopsys translate_off
	`endif
                          ,
                          .clkswitch(1'b0),
                          .configupdate(1'b0),
                          .pfdena(1'b1),
                          .phasecounterselect({3{1'b0}}),
                          .phasestep(1'b0),
                          .phaseupdown(1'b0),
                          .scanclk(1'b0),
                          .scanclkena(1'b1),
                          .scandata(1'b0)
	`ifndef FORMAL_VERIFICATION
                          // synopsys translate_on
	`endif
                      );
    defparam
        pll7.bandwidth_type = "auto",
        pll7.clk0_divide_by = 1,
        pll7.clk0_duty_cycle = 50,
        pll7.clk0_multiply_by = 1,
        pll7.clk0_phase_shift = "0",
        pll7.clk1_divide_by = 25,
        pll7.clk1_duty_cycle = 50,
        pll7.clk1_multiply_by = 1,
        pll7.clk1_phase_shift = "0",
        pll7.compensate_clock = "clk0",
        pll7.inclk0_input_frequency = 20000,
        pll7.operation_mode = "normal",
        pll7.pll_type = "auto",
        pll7.lpm_type = "fiftyfivenm_pll";
    assign
        clk = {wire_pll7_clk[4:0]},
        locked = (wire_pll7_locked & pll_lock_sync);
endmodule //adc_altpll_0_altpll_nc92

module  adc_altpll_0
    (
        address,
        areset,
        c0,
        c1,
        clk,
        locked,
        phasecounterselect,
        phasedone,
        phasestep,
        phaseupdown,
        read,
        readdata,
        reset,
        scanclk,
        write,
        writedata) /* synthesis synthesis_clearbox=1 */;
    input   [1:0]  address;
    input   areset;
    output   c0;
    output   c1;
    input   clk;
    output   locked;
    input   [2:0]  phasecounterselect;
    output   phasedone;
    input   phasestep;
    input   phaseupdown;
    input   read;
    output   [31:0]  readdata;
    input   reset;
    input   scanclk;
    input   write;
    input   [31:0]  writedata;

    wire  wire_stdsync2_dout;
    wire  [4:0]   wire_sd1_clk;
    wire  wire_sd1_locked;
    (* ALTERA_ATTRIBUTE = {"POWER_UP_LEVEL=HIGH"} *)
    reg	pfdena_reg;
    wire	wire_pfdena_reg_ena;
    reg	prev_reset;
    wire  w_locked;
    wire  w_pfdena;
    wire  w_phasedone;
    wire  w_pll_areset_in;
    wire  w_reset;
    wire  w_select_control;
    wire  w_select_status;

    adc_altpll_0_stdsync_sv6   stdsync2
                               (
                                   .clk(clk),
                                   .din(wire_sd1_locked),
                                   .dout(wire_stdsync2_dout),
                                   .reset_n((~ reset)));
    adc_altpll_0_altpll_nc92   sd1
                               (
                                   .areset((w_pll_areset_in | areset)),
                                   .clk(wire_sd1_clk),
                                   .inclk({{1{1'b0}}, clk}),
                                   .locked(wire_sd1_locked));
    // synopsys translate_off
    initial
        pfdena_reg = {1{1'b1}};
    // synopsys translate_on
    always @ ( posedge clk or  posedge reset)
        if (reset == 1'b1) pfdena_reg <= {1{1'b1}};
        else if  (wire_pfdena_reg_ena == 1'b1)   pfdena_reg <= writedata[1];
    assign
        wire_pfdena_reg_ena = (write & w_select_control);
    // synopsys translate_off
    initial
        prev_reset = 0;
    // synopsys translate_on
    always @ ( posedge clk or  posedge reset)
        if (reset == 1'b1) prev_reset <= 1'b0;
        else  prev_reset <= w_reset;
    assign
        c0 = wire_sd1_clk[0],
        c1 = wire_sd1_clk[1],
        locked = wire_sd1_locked,
        phasedone = 1'b0,
        readdata = {{30{1'b0}}, (read & ((w_select_control & w_pfdena) | (w_select_status & w_phasedone))), (read & ((w_select_control & w_pll_areset_in) | (w_select_status & w_locked)))},
        w_locked = wire_stdsync2_dout,
        w_pfdena = pfdena_reg,
        w_phasedone = 1'b1,
        w_pll_areset_in = prev_reset,
        w_reset = ((write & w_select_control) & writedata[0]),
        w_select_control = ((~ address[1]) & address[0]),
        w_select_status = ((~ address[1]) & (~ address[0]));
endmodule //adc_altpll_0


module adc_modular_adc_0 #(
        parameter is_this_first_or_second_adc = 1
    ) (
        input  wire        clock_clk,              //          clock.clk
        input  wire        reset_sink_reset_n,     //     reset_sink.reset_n
        input  wire        adc_pll_clock_clk,      //  adc_pll_clock.clk
        input  wire        adc_pll_locked_export,  // adc_pll_locked.export
        input  wire        command_valid,          //        command.valid
        input  wire [4:0]  command_channel,        //               .channel
        input  wire        command_startofpacket,  //               .startofpacket
        input  wire        command_endofpacket,    //               .endofpacket
        output wire        command_ready,          //               .ready
        output wire        response_valid,         //       response.valid
        output wire [4:0]  response_channel,       //               .channel
        output wire [11:0] response_data,          //               .data
        output wire        response_startofpacket, //               .startofpacket
        output wire        response_endofpacket    //               .endofpacket
    );

    generate
        if (is_this_first_or_second_adc != 1)
        begin
            initial begin
                $display("Generated module instantiated with wrong parameters");
                $stop;
            end
            instantiated_with_wrong_parameters_error_see_comment_above
                is_this_first_or_second_adc_check ( .error(1'b1) );
        end
    endgenerate

    altera_modular_adc_control #(
                                   .clkdiv                          (4),
                                   .tsclkdiv                        (0),
                                   .tsclksel                        (1),
                                   .hard_pwd                        (0),
                                   .prescalar                       (0),
                                   .refsel                          (0),
                                   .device_partname_fivechar_prefix ("10M50"),
                                   .is_this_first_or_second_adc     (1),
                                   .analog_input_pin_mask           (65536),
                                   .dual_adc_mode                   (0),
                                   .enable_usr_sim                  (0),
                                   .reference_voltage_sim           (49648),
                                   .simfilename_ch0                 (""),
                                   .simfilename_ch1                 (""),
                                   .simfilename_ch2                 (""),
                                   .simfilename_ch3                 (""),
                                   .simfilename_ch4                 (""),
                                   .simfilename_ch5                 (""),
                                   .simfilename_ch6                 (""),
                                   .simfilename_ch7                 (""),
                                   .simfilename_ch8                 (""),
                                   .simfilename_ch9                 (""),
                                   .simfilename_ch10                (""),
                                   .simfilename_ch11                (""),
                                   .simfilename_ch12                (""),
                                   .simfilename_ch13                (""),
                                   .simfilename_ch14                (""),
                                   .simfilename_ch15                (""),
                                   .simfilename_ch16                ("")
                               ) control_internal (
                                   .clk               (clock_clk),              //         clock.clk
                                   .cmd_valid         (command_valid),          //       command.valid
                                   .cmd_channel       (command_channel),        //              .channel
                                   .cmd_sop           (command_startofpacket),  //              .startofpacket
                                   .cmd_eop           (command_endofpacket),    //              .endofpacket
                                   .cmd_ready         (command_ready),          //              .ready
                                   .rst_n             (reset_sink_reset_n),     //    reset_sink.reset_n
                                   .rsp_valid         (response_valid),         //      response.valid
                                   .rsp_channel       (response_channel),       //              .channel
                                   .rsp_data          (response_data),          //              .data
                                   .rsp_sop           (response_startofpacket), //              .startofpacket
                                   .rsp_eop           (response_endofpacket),   //              .endofpacket
                                   .clk_in_pll_c0     (adc_pll_clock_clk),      // adc_pll_clock.clk
                                   .clk_in_pll_locked (adc_pll_locked_export),  //   conduit_end.export
                                   .sync_valid        (),                       //   (terminated)
                                   .sync_ready        (1'b0)                    //   (terminated)
                               );

endmodule

module altera_modular_adc_control #(
        parameter clkdiv        = 1,
        parameter tsclkdiv      = 0,
        parameter tsclksel      = 0,
        parameter prescalar     = 0,
        parameter refsel        = 0,
        parameter device_partname_fivechar_prefix   = "10M08",
        parameter is_this_first_or_second_adc = 1,
        parameter analog_input_pin_mask = 17'h0,
        parameter hard_pwd = 0,
        parameter dual_adc_mode = 0,
        parameter enable_usr_sim = 0,
        parameter reference_voltage_sim = 65536,
        parameter simfilename_ch0 = "simfilename_ch0",
        parameter simfilename_ch1 = "simfilename_ch1",
        parameter simfilename_ch2 = "simfilename_ch2",
        parameter simfilename_ch3 = "simfilename_ch3",
        parameter simfilename_ch4 = "simfilename_ch4",
        parameter simfilename_ch5 = "simfilename_ch5",
        parameter simfilename_ch6 = "simfilename_ch6",
        parameter simfilename_ch7 = "simfilename_ch7",
        parameter simfilename_ch8 = "simfilename_ch8",
        parameter simfilename_ch9 = "simfilename_ch9",
        parameter simfilename_ch10 = "simfilename_ch10",
        parameter simfilename_ch11 = "simfilename_ch11",
        parameter simfilename_ch12 = "simfilename_ch12",
        parameter simfilename_ch13 = "simfilename_ch13",
        parameter simfilename_ch14 = "simfilename_ch14",
        parameter simfilename_ch15 = "simfilename_ch15",
        parameter simfilename_ch16 = "simfilename_ch16"
    ) (
        input           clk,
        input           rst_n,
        input           clk_in_pll_c0,
        input           clk_in_pll_locked,
        input           cmd_valid,
        input [4:0]     cmd_channel,
        input           cmd_sop,
        input           cmd_eop,
        input           sync_ready,

        output          cmd_ready,
        output          rsp_valid,
        output [4:0]    rsp_channel,
        output [11:0]   rsp_data,
        output          rsp_sop,
        output          rsp_eop,
        output          sync_valid

    );

    wire        clkout_adccore;
    wire        eoc;
    wire [11:0] dout;
    wire [4:0]  chsel;
    wire        soc;
    wire        tsen;
    wire        usr_pwd;

    altera_modular_adc_control_fsm #(
                                       .is_this_first_or_second_adc    (is_this_first_or_second_adc),
                                       .dual_adc_mode                  (dual_adc_mode)
                                   ) u_control_fsm (
                                       // inputs
                                       .clk                (clk),
                                       .rst_n              (rst_n),
                                       .clk_in_pll_locked  (clk_in_pll_locked),
                                       .cmd_valid          (cmd_valid),
                                       .cmd_channel        (cmd_channel),
                                       .cmd_sop            (cmd_sop),
                                       .cmd_eop            (cmd_eop),
                                       .clk_dft            (clkout_adccore),
                                       .eoc                (eoc),
                                       .dout               (dout),
                                       .sync_ready         (sync_ready),
                                       // outputs
                                       .rsp_valid          (rsp_valid),
                                       .rsp_channel        (rsp_channel),
                                       .rsp_data           (rsp_data),
                                       .rsp_sop            (rsp_sop),
                                       .rsp_eop            (rsp_eop),
                                       .cmd_ready          (cmd_ready),
                                       .chsel              (chsel),
                                       .soc                (soc),
                                       .usr_pwd            (usr_pwd),
                                       .tsen               (tsen),
                                       .sync_valid         (sync_valid)
                                   );


    fiftyfivenm_adcblock_top_wrapper #(
                                         .device_partname_fivechar_prefix (device_partname_fivechar_prefix),
                                         .clkdiv                          (clkdiv),
                                         .tsclkdiv                        (tsclkdiv),
                                         .tsclksel                        (tsclksel),
                                         .refsel                          (refsel),
                                         .prescalar                       (prescalar),
                                         .is_this_first_or_second_adc     (is_this_first_or_second_adc),
                                         .analog_input_pin_mask           (analog_input_pin_mask),
                                         .hard_pwd                        (hard_pwd),
                                         .enable_usr_sim                  (enable_usr_sim),
                                         .reference_voltage_sim           (reference_voltage_sim),
                                         .simfilename_ch0                 (simfilename_ch0),
                                         .simfilename_ch1                 (simfilename_ch1),
                                         .simfilename_ch2                 (simfilename_ch2),
                                         .simfilename_ch3                 (simfilename_ch3),
                                         .simfilename_ch4                 (simfilename_ch4),
                                         .simfilename_ch5                 (simfilename_ch5),
                                         .simfilename_ch6                 (simfilename_ch6),
                                         .simfilename_ch7                 (simfilename_ch7),
                                         .simfilename_ch8                 (simfilename_ch8),
                                         .simfilename_ch9                 (simfilename_ch9),
                                         .simfilename_ch10                (simfilename_ch10),
                                         .simfilename_ch11                (simfilename_ch11),
                                         .simfilename_ch12                (simfilename_ch12),
                                         .simfilename_ch13                (simfilename_ch13),
                                         .simfilename_ch14                (simfilename_ch14),
                                         .simfilename_ch15                (simfilename_ch15),
                                         .simfilename_ch16                (simfilename_ch16)
                                     ) adc_inst (
                                         //.reset              (reset),
                                         .chsel              (chsel),                        // 5-bits channel selection.
                                         .soc                (soc),                          // signal Start-of-Conversion to ADC
                                         .eoc                (eoc),                          // signal end of conversion. Data can be latched on the positive edge of clkout_adccore after this signal becomes high.  EOC becomes low at every positive edge of the clkout_adccore signal.
                                         .dout               (dout),                         // 12-bits DOUT valid after EOC rise, still valid at falling edge, but not before the next EOC rising edge
                                         .usr_pwd            (usr_pwd),                      // User Power Down during run time.  0 = Power Up;  1 = Power Down.
                                         .tsen               (tsen),                         // MUST power down ADC before changing TSEN.  0 = Normal Mode; 1 = Temperature Sensing Mode.
                                         .clkout_adccore     (clkout_adccore),               // Output clock from the clock divider
                                         .clkin_from_pll_c0  (clk_in_pll_c0)               // Clock source from PLL1/3 c-counter[0]
                                         //.dout_ch            (dout_ch)                     // Indicate dout is for which chsel
                                     );

endmodule



module altera_modular_adc_control_fsm #(
        parameter is_this_first_or_second_adc = 1,
        parameter dual_adc_mode = 0
    ) (
        input               clk,
        input               rst_n,
        input               clk_in_pll_locked,
        input               cmd_valid,
        input [4:0]         cmd_channel,
        input               cmd_sop,
        input               cmd_eop,
        input               clk_dft,
        input               eoc,
        input [11:0]        dout,
        input               sync_ready,

        output reg          rsp_valid,
        output reg [4:0]    rsp_channel,
        output reg [11:0]   rsp_data,
        output reg          rsp_sop,
        output reg          rsp_eop,
        output reg          cmd_ready,
        output reg [4:0]    chsel,
        output reg          soc,
        output reg          usr_pwd,
        output reg          tsen,
        output reg          sync_valid

    );

    reg [4:0]   ctrl_state;
    reg [4:0]   ctrl_state_nxt;
    reg         clk_dft_synch_dly;
    reg         eoc_synch_dly;
    reg [4:0]   chsel_nxt;
    reg         soc_nxt;
    reg         usr_pwd_nxt;
    reg         tsen_nxt;
    reg         prev_cmd_is_ts;
    reg         cmd_fetched;
    reg         pend;
    reg [4:0]   cmd_channel_dly;
    reg         cmd_sop_dly;
    reg         cmd_eop_dly;
    reg [7:0]   int_timer;
    reg [17:0]  avrg_sum;
    reg         avrg_cnt_done;
    reg         frst_64_ptr_done;
    reg         conv_dly1_s_flp;
    reg [11:0]  dout_flp;
    reg [4:0]   prev_ctrl_state;
    reg [4:0]   sync_ctrl_state;
    reg [4:0]   sync_ctrl_state_nxt;

    wire        clk_dft_synch;
    wire        eoc_synch;
    wire        clk_dft_lh;
    wire        clk_dft_hl;
    wire        eoc_hl;
    wire        cmd_is_rclb;
    wire        cmd_is_ts;
    wire        arc_conv_conv_dly1;
    wire        arc_sync1_conv_dly1;
    wire        arc_wait_pend_wait_pend_dly1;
    wire        arc_sync1_wait_pend_dly1;
    wire        arc_to_conv;
    wire        arc_to_avrg_cnt;
    wire        load_rsp;
    wire        load_cmd_ready;
    wire        arc_getcmd_w_pwrdwn;
    wire        arc_getcmd_pwrdwn;
    wire        load_cmd_fetched;
    wire        load_int_timer;
    wire        incr_int_timer;
    wire        arc_out_from_pwrup_soc;
    wire        clr_cmd_fetched;
    wire        adc_change_mode;
    wire        add_avrg_sum;
    wire        add_avrg_sum_run;
    wire        clear_avrg_sum;
    wire        clear_avrg_cnt_done;
    wire        set_frst_64_ptr_done;
    wire        clear_frst_64_ptr_done;
    wire [11:0] fifo_q;
    wire        fifo_sclr;
    wire        fifo_rdreq;
    wire        fifo_wrreq;
    wire        putresp_s;
    wire        putresp_pend_s;
    wire        pwrdwn_s;
    wire        pwrdwn_tsen_s;
    wire        avrg_cnt_s;
    wire        wait_pend_dly1_s;
    wire        conv_dly1_s;
    wire        conv_s;
    wire        putresp_dly3_s;
    wire        load_dout;
    wire        avrg_enable;
    wire [11:0] rsp_data_nxt;

    localparam [4:0]    IDLE                = 5'b00000;
    localparam [4:0]    PWRDWN              = 5'b00001;
    localparam [4:0]    PWRDWN_TSEN         = 5'b00010;
    localparam [4:0]    PWRDWN_DONE         = 5'b00011;
    localparam [4:0]    PWRUP_CH            = 5'b00100;
    localparam [4:0]    PWRUP_SOC           = 5'b00101;
    localparam [4:0]    WAIT                = 5'b00110;
    localparam [4:0]    GETCMD              = 5'b00111;
    localparam [4:0]    GETCMD_W            = 5'b01000;
    localparam [4:0]    PRE_CONV            = 5'b01001;
    localparam [4:0]    CONV                = 5'b01010; // Drive chsel. Get out of this state when falling edge of EOC detected (DOUT is ready for sample)
    // Read averaging fifo.
    // Capture DOUT into dout internal buffer register (dout_flp)
    localparam [4:0]    CONV_DLY1           = 5'b01011; // Additional state for processing when DOUT is ready. Perform averaging calculation (adds and minus operation).
    localparam [4:0]    PUTRESP             = 5'b01100; // Load response
    localparam [4:0]    PUTRESP_DLY1        = 5'b01101;
    localparam [4:0]    PUTRESP_DLY2        = 5'b01110;
    localparam [4:0]    PUTRESP_DLY3        = 5'b01111;
    localparam [4:0]    WAIT_PEND           = 5'b10000; // Get out of this state when falling edge of EOC detected (DOUT is ready for sample)
    // Read averaging fifo.
    // Capture DOUT into dout internal buffer register (dout_flp)
    localparam [4:0]    WAIT_PEND_DLY1      = 5'b10001; // Additional state for processing when DOUT is ready. Perform averaging calculation (adds and minus operation).
    localparam [4:0]    PUTRESP_PEND        = 5'b10010; // Load response
    localparam [4:0]    AVRG_CNT            = 5'b10011;
    localparam [4:0]    SYNC1               = 5'b10100; // Allocates 1 soft ip clock mismatch due to asynchronous between soft ip clock and ADC clock domain

    localparam [7:0]    NUM_AVRG_POINTS     = 8'd64;

    //--------------------------------------------------------------------------------------------//
    // Double Synchronize control signal from ADC hardblock
    //--------------------------------------------------------------------------------------------//
    altera_std_synchronizer #(
                                .depth    (2)
                            ) u_clk_dft_synchronizer (
                                .clk        (clk),
                                .reset_n    (rst_n),
                                .din        (clk_dft),
                                .dout       (clk_dft_synch)
                            );

    altera_std_synchronizer #(
                                .depth    (2)
                            ) u_eoc_synchronizer (
                                .clk        (clk),
                                .reset_n    (rst_n),
                                .din        (eoc),
                                .dout       (eoc_synch)
                            );



    //--------------------------------------------------------------------------------------------//
    // Edge detection for both synchronized clk_dft and eoc
    //--------------------------------------------------------------------------------------------//
    always @(posedge clk or negedge rst_n) begin
        if (!rst_n) begin
            clk_dft_synch_dly   <= 1'b0;
            eoc_synch_dly       <= 1'b0;
        end
        else begin
            clk_dft_synch_dly   <= clk_dft_synch;
            eoc_synch_dly       <= eoc_synch;
        end
    end

    assign clk_dft_lh   = clk_dft_synch & ~clk_dft_synch_dly;
    assign clk_dft_hl   = ~clk_dft_synch & clk_dft_synch_dly;
    assign eoc_hl       = ~eoc_synch & eoc_synch_dly;


    //--------------------------------------------------------------------------------------------//
    // Dual ADC
    //--------------------------------------------------------------------------------------------//

    generate
        if (dual_adc_mode == 1) begin

            // Buffer up ctrl_state
            // To be used when both ADC is out of sync
            always @(posedge clk or negedge rst_n) begin
                if (!rst_n)
                    prev_ctrl_state   <= IDLE;
                else
                    prev_ctrl_state   <= ctrl_state;
            end

            // Buffer up ctrl_state
            // To be used when both ADC mismatches by 1 soft ip clock
            always @(posedge clk or negedge rst_n) begin
                if (!rst_n)
                    sync_ctrl_state   <= IDLE;
                else
                    sync_ctrl_state   <= sync_ctrl_state_nxt;
            end

        end
        else begin

            always @* begin
                prev_ctrl_state = 5'h0;
                sync_ctrl_state = 5'h0;
            end

        end
    endgenerate



    //--------------------------------------------------------------------------------------------//
    // Main FSM
    //--------------------------------------------------------------------------------------------//
    always @(posedge clk or negedge rst_n) begin
        if (!rst_n)
            ctrl_state   <= IDLE;
        else
            ctrl_state   <= ctrl_state_nxt;
    end


    always @* begin

        // Default assignment, perform assignment only at relevant state
        sync_ctrl_state_nxt = sync_ctrl_state;
        sync_valid          = 1'b0;

        case (ctrl_state)
            IDLE: begin
                if (clk_in_pll_locked)
                    ctrl_state_nxt = PWRDWN;
                else
                    ctrl_state_nxt = IDLE;
            end

            PWRDWN: begin
                if (int_timer[6])
                    ctrl_state_nxt = PWRDWN_TSEN;
                else
                    ctrl_state_nxt = PWRDWN;
            end

            PWRDWN_TSEN: begin
                if (int_timer[7])
                    ctrl_state_nxt = PWRDWN_DONE;
                else
                    ctrl_state_nxt = PWRDWN_TSEN;
            end

            PWRDWN_DONE: begin
                if (dual_adc_mode == 1) begin
                    if (clk_dft_lh) begin
                        if (sync_ready)
                            ctrl_state_nxt = PWRUP_CH;
                        else
                            ctrl_state_nxt = SYNC1;
                    end
                    else begin
                        ctrl_state_nxt = PWRDWN_DONE;
                    end

                    if (clk_dft_lh) begin
                        sync_ctrl_state_nxt = PWRUP_CH;
                        sync_valid          = 1'b1;
                    end

                end
                else begin
                    if (clk_dft_lh)
                        ctrl_state_nxt = PWRUP_CH;
                    else
                        ctrl_state_nxt = PWRDWN_DONE;
                end
            end

            PWRUP_CH: begin
                if (dual_adc_mode == 1) begin
                    if (clk_dft_hl) begin
                        if (sync_ready)
                            ctrl_state_nxt = PWRUP_SOC;
                        else
                            ctrl_state_nxt = SYNC1;
                    end
                    else begin
                        ctrl_state_nxt = PWRUP_CH;
                    end

                    if (clk_dft_hl) begin
                        sync_ctrl_state_nxt = PWRUP_SOC;
                        sync_valid          = 1'b1;
                    end

                end
                else begin
                    if (clk_dft_hl)
                        ctrl_state_nxt = PWRUP_SOC;
                    else
                        ctrl_state_nxt = PWRUP_CH;
                end
            end

            PWRUP_SOC: begin
                if (dual_adc_mode == 1) begin
                    if (eoc_hl) begin
                        if (sync_ready) begin
                            if (cmd_fetched & ~cmd_is_rclb)
                                ctrl_state_nxt = CONV;
                            else if (cmd_fetched & cmd_is_rclb)
                                ctrl_state_nxt = PUTRESP;
                            else if (cmd_valid)
                                ctrl_state_nxt = GETCMD;
                            else
                                ctrl_state_nxt = WAIT;
                        end
                        else begin
                            ctrl_state_nxt = SYNC1;
                        end
                    end
                    else begin
                        ctrl_state_nxt = PWRUP_SOC;
                    end

                    if (eoc_hl) begin
                        if (cmd_fetched & ~cmd_is_rclb)
                            sync_ctrl_state_nxt = CONV;
                        else if (cmd_fetched & cmd_is_rclb)
                            sync_ctrl_state_nxt = PUTRESP;
                        else if (cmd_valid)
                            sync_ctrl_state_nxt = GETCMD;
                        else
                            sync_ctrl_state_nxt = WAIT;

                        sync_valid  = 1'b1;
                    end

                end
                else begin
                    if (cmd_fetched & ~cmd_is_rclb & eoc_hl)
                        ctrl_state_nxt = CONV;
                    else if (cmd_fetched & cmd_is_rclb & eoc_hl)
                        ctrl_state_nxt = PUTRESP;
                    else if (cmd_valid & eoc_hl)
                        ctrl_state_nxt = GETCMD;
                    else if (eoc_hl)
                        ctrl_state_nxt = WAIT;
                    else
                        ctrl_state_nxt = PWRUP_SOC;
                end
            end

            SYNC1: begin
                if (sync_ready)
                    ctrl_state_nxt = sync_ctrl_state;   // mismatches by 1 soft ip clock, proceed to next state
                else
                    ctrl_state_nxt = prev_ctrl_state;   // Both ADC is out of sync, go back to previous state

                sync_valid  = 1'b1;

            end

            WAIT: begin
                if (cmd_valid)
                    ctrl_state_nxt = GETCMD_W;
                else
                    ctrl_state_nxt = WAIT;
            end

            GETCMD_W: begin
                if (cmd_is_rclb | adc_change_mode)
                    ctrl_state_nxt = PWRDWN;
                else
                    ctrl_state_nxt = PRE_CONV;
            end

            PRE_CONV: begin
                if (dual_adc_mode == 1) begin
                    if (eoc_hl) begin
                        if (sync_ready)
                            ctrl_state_nxt = CONV;
                        else
                            ctrl_state_nxt = SYNC1;
                    end
                    else begin
                        ctrl_state_nxt = PRE_CONV;
                    end

                    if (eoc_hl) begin
                        sync_ctrl_state_nxt = CONV;
                        sync_valid          = 1'b1;
                    end

                end
                else begin
                    if (eoc_hl)
                        ctrl_state_nxt = CONV;
                    else
                        ctrl_state_nxt = PRE_CONV;
                end
            end

            GETCMD: begin
                if ((cmd_is_rclb | adc_change_mode) & ~pend)
                    ctrl_state_nxt = PWRDWN;
                else if ((cmd_is_rclb | adc_change_mode) & pend)
                    ctrl_state_nxt = WAIT_PEND;
                else
                    ctrl_state_nxt = CONV;
            end

            CONV: begin
                if (dual_adc_mode == 1) begin
                    if (eoc_hl) begin
                        if (sync_ready) begin
                            if (avrg_enable & ~avrg_cnt_done)
                                ctrl_state_nxt = AVRG_CNT;
                            else
                                ctrl_state_nxt = CONV_DLY1;
                        end
                        else begin
                            ctrl_state_nxt = SYNC1;
                        end
                    end
                    else begin
                        ctrl_state_nxt = CONV;
                    end

                    if (eoc_hl) begin
                        if (avrg_enable & ~avrg_cnt_done)
                            sync_ctrl_state_nxt = AVRG_CNT;
                        else
                            sync_ctrl_state_nxt = CONV_DLY1;

                        sync_valid  = 1'b1;
                    end

                end
                else begin
                    if (eoc_hl & avrg_enable & ~avrg_cnt_done)
                        ctrl_state_nxt = AVRG_CNT;
                    else if (eoc_hl)
                        ctrl_state_nxt = CONV_DLY1;
                    else
                        ctrl_state_nxt = CONV;
                end
            end

            AVRG_CNT: begin
                ctrl_state_nxt = CONV;
            end

            CONV_DLY1: begin
                ctrl_state_nxt = PUTRESP;
            end

            PUTRESP: begin
                ctrl_state_nxt = PUTRESP_DLY1;
            end

            PUTRESP_DLY1: begin
                ctrl_state_nxt = PUTRESP_DLY2;
            end

            PUTRESP_DLY2: begin
                ctrl_state_nxt = PUTRESP_DLY3;
            end

            PUTRESP_DLY3: begin
                if (cmd_valid)
                    ctrl_state_nxt = GETCMD;
                else if (pend)
                    ctrl_state_nxt = WAIT_PEND;
                else
                    ctrl_state_nxt = WAIT;
            end

            WAIT_PEND: begin
                if (dual_adc_mode == 1) begin
                    if (eoc_hl) begin
                        if (sync_ready)
                            ctrl_state_nxt = WAIT_PEND_DLY1;
                        else
                            ctrl_state_nxt = SYNC1;
                    end
                    else begin
                        ctrl_state_nxt = WAIT_PEND;
                    end

                    if (eoc_hl) begin
                        sync_ctrl_state_nxt = WAIT_PEND_DLY1;
                        sync_valid          = 1'b1;
                    end

                end
                else begin
                    if (eoc_hl)
                        ctrl_state_nxt = WAIT_PEND_DLY1;
                    else
                        ctrl_state_nxt = WAIT_PEND;
                end
            end

            WAIT_PEND_DLY1: begin
                ctrl_state_nxt = PUTRESP_PEND;
            end

            PUTRESP_PEND: begin
                if (cmd_valid)
                    ctrl_state_nxt = GETCMD;
                else
                    ctrl_state_nxt = WAIT;
            end

            default: begin
                ctrl_state_nxt = IDLE;
            end

        endcase
    end



    always @* begin
        chsel_nxt       = chsel;
        soc_nxt         = soc;
        usr_pwd_nxt     = usr_pwd;
        tsen_nxt        = tsen;

        case (ctrl_state_nxt)
            IDLE: begin
                chsel_nxt   = 5'b11110;
                soc_nxt     = 1'b0;
                usr_pwd_nxt = 1'b1;
                tsen_nxt    = 1'b0;
            end

            PWRDWN: begin
                chsel_nxt   = chsel;
                soc_nxt     = 1'b0;
                usr_pwd_nxt = 1'b1;
                tsen_nxt    = tsen;
            end

            PWRDWN_TSEN: begin
                chsel_nxt   = chsel;
                soc_nxt     = 1'b0;
                usr_pwd_nxt = 1'b1;
                if (cmd_fetched & cmd_is_ts)        // Transition to TS mode
                    tsen_nxt    = 1'b1;
                else if (cmd_fetched & cmd_is_rclb) // In recalibration mode, maintain previous TSEN setting
                    tsen_nxt    = tsen;
                else
                    tsen_nxt    = 1'b0;             // Transition to Normal mode
            end

            PWRDWN_DONE: begin
                chsel_nxt   = chsel;
                soc_nxt     = 1'b0;
                usr_pwd_nxt = 1'b0;
                tsen_nxt    = tsen;
            end

            PWRUP_CH: begin
                chsel_nxt   = 5'b11110;
                soc_nxt     = soc;
                usr_pwd_nxt = 1'b0;
                tsen_nxt    = tsen;
            end

            PWRUP_SOC: begin
                chsel_nxt   = chsel;
                soc_nxt     = 1'b1;
                usr_pwd_nxt = usr_pwd;
                tsen_nxt    = tsen;
            end

            SYNC1: begin
                chsel_nxt   = chsel;
                soc_nxt     = soc;
                usr_pwd_nxt = usr_pwd;
                tsen_nxt    = tsen;
            end

            WAIT: begin
                chsel_nxt   = chsel;
                soc_nxt     = soc;
                usr_pwd_nxt = usr_pwd;
                tsen_nxt    = tsen;
            end

            GETCMD_W: begin
                chsel_nxt   = chsel;
                soc_nxt     = soc;
                usr_pwd_nxt = usr_pwd;
                tsen_nxt    = tsen;
            end

            PRE_CONV: begin
                chsel_nxt   = chsel;
                soc_nxt     = soc;
                usr_pwd_nxt = usr_pwd;
                tsen_nxt    = tsen;
            end

            GETCMD: begin
                chsel_nxt   = chsel;
                soc_nxt     = soc;
                usr_pwd_nxt = usr_pwd;
                tsen_nxt    = tsen;
            end

            CONV: begin
                chsel_nxt   = cmd_channel;
                soc_nxt     = soc;
                usr_pwd_nxt = usr_pwd;
                tsen_nxt    = tsen;
            end

            AVRG_CNT: begin
                chsel_nxt   = cmd_channel;
                soc_nxt     = soc;
                usr_pwd_nxt = usr_pwd;
                tsen_nxt    = tsen;
            end

            CONV_DLY1: begin
                chsel_nxt   = cmd_channel;
                soc_nxt     = soc;
                usr_pwd_nxt = usr_pwd;
                tsen_nxt    = tsen;
            end

            PUTRESP: begin
                chsel_nxt   = chsel;
                soc_nxt     = soc;
                usr_pwd_nxt = usr_pwd;
                tsen_nxt    = tsen;
            end

            PUTRESP_DLY1: begin
                chsel_nxt   = chsel;
                soc_nxt     = soc;
                usr_pwd_nxt = usr_pwd;
                tsen_nxt    = tsen;
            end

            PUTRESP_DLY2: begin
                chsel_nxt   = chsel;
                soc_nxt     = soc;
                usr_pwd_nxt = usr_pwd;
                tsen_nxt    = tsen;
            end

            PUTRESP_DLY3: begin
                chsel_nxt   = chsel;
                soc_nxt     = soc;
                usr_pwd_nxt = usr_pwd;
                tsen_nxt    = tsen;
            end

            WAIT_PEND: begin
                //chsel_nxt   = chsel;
                chsel_nxt   = 5'b11110; // The reason for this change is to support ADC's simulation model (case:226093).
                // During the final sampling cycle which meant to complete the pending ADC sampling (ADC output is one cycle delay in nature),
                // we assign a dummy channel value instead of maintaining the previous channel value. Functionally, it does not matter.
                // But it does matter to simulation model where it keep popping up the expected value from user's simulation file based on current channel value.
                // This will avoid the simulation model from incorrectly popping out the value from previous channel twice during ADC mode transition.
                soc_nxt     = soc;
                usr_pwd_nxt = usr_pwd;
                tsen_nxt    = tsen;
            end

            WAIT_PEND_DLY1: begin
                chsel_nxt   = chsel;
                soc_nxt     = soc;
                usr_pwd_nxt = usr_pwd;
                tsen_nxt    = tsen;
            end

            PUTRESP_PEND: begin
                chsel_nxt   = chsel;
                soc_nxt     = soc;
                usr_pwd_nxt = usr_pwd;
                tsen_nxt    = tsen;
            end

            default: begin
                chsel_nxt   = 5'bx;
                soc_nxt     = 1'bx;
                usr_pwd_nxt = 1'bx;
                tsen_nxt    = 1'bx;
            end

        endcase
    end



    always @(posedge clk or negedge rst_n) begin
        if (!rst_n) begin
            chsel       <= 5'b11110;
            soc         <= 1'b0;
            usr_pwd     <= 1'b1;
            tsen        <= 1'b0;
        end
        else begin
            chsel       <= chsel_nxt;
            soc         <= soc_nxt;
            usr_pwd     <= usr_pwd_nxt;
            tsen        <= tsen_nxt;

        end
    end



    assign arc_conv_conv_dly1               = (ctrl_state == CONV) & (ctrl_state_nxt == CONV_DLY1);
    assign arc_wait_pend_wait_pend_dly1     = (ctrl_state == WAIT_PEND) & (ctrl_state_nxt == WAIT_PEND_DLY1);
    assign arc_to_avrg_cnt                  = ((ctrl_state == CONV) & (ctrl_state_nxt == AVRG_CNT)) | ((ctrl_state == SYNC1) & (ctrl_state_nxt == AVRG_CNT));

    assign arc_sync1_conv_dly1              = (ctrl_state == SYNC1) & (ctrl_state_nxt == CONV_DLY1);        // prev_ctrl_state is guaranteed by design to be CONV
    assign arc_sync1_wait_pend_dly1         = (ctrl_state == SYNC1) & (ctrl_state_nxt == WAIT_PEND_DLY1);   // prev_ctrl_state is guaranteed by design to be WAIT_PEND


    assign putresp_s        = (ctrl_state == PUTRESP);
    assign putresp_pend_s   = (ctrl_state == PUTRESP_PEND);
    assign pwrdwn_s         = (ctrl_state == PWRDWN);
    assign pwrdwn_tsen_s    = (ctrl_state == PWRDWN_TSEN);
    assign avrg_cnt_s       = (ctrl_state == AVRG_CNT);
    assign wait_pend_dly1_s = (ctrl_state == WAIT_PEND_DLY1);
    assign conv_dly1_s      = (ctrl_state == CONV_DLY1);
    assign conv_s           = (ctrl_state == CONV);
    assign putresp_dly3_s   = (ctrl_state == PUTRESP_DLY3);



    assign load_rsp                     = (putresp_s & ~cmd_is_rclb & pend) | putresp_pend_s;
    assign load_dout                    = ((arc_conv_conv_dly1 | arc_sync1_conv_dly1) & ~cmd_is_rclb & pend) | arc_wait_pend_wait_pend_dly1 | arc_sync1_wait_pend_dly1 | ((int_timer != 8'h0) & arc_to_avrg_cnt);
    assign load_cmd_ready               = putresp_s;
    assign arc_to_conv                  = (ctrl_state != CONV) & (ctrl_state != AVRG_CNT) & ~((ctrl_state == SYNC1) & (prev_ctrl_state == CONV)) & (ctrl_state_nxt == CONV);

    assign arc_getcmd_w_pwrdwn          = (ctrl_state == GETCMD_W) & (ctrl_state_nxt == PWRDWN);
    assign arc_getcmd_pwrdwn            = (ctrl_state == GETCMD) & (ctrl_state_nxt == PWRDWN);
    assign load_cmd_fetched             = arc_getcmd_w_pwrdwn | arc_getcmd_pwrdwn;
    assign load_int_timer               = arc_getcmd_w_pwrdwn | arc_getcmd_pwrdwn | arc_to_conv; // arc_to_conv is added for averaging
    assign incr_int_timer               = pwrdwn_s | pwrdwn_tsen_s | avrg_cnt_s;

    assign arc_out_from_pwrup_soc       = ((ctrl_state == PWRUP_SOC) & (ctrl_state_nxt != PWRUP_SOC) & (ctrl_state_nxt != SYNC1)) |
           ((ctrl_state == SYNC1) & (prev_ctrl_state == PWRUP_SOC) & (ctrl_state_nxt != PWRUP_SOC));
    assign clr_cmd_fetched              = arc_out_from_pwrup_soc;

    assign cmd_is_rclb      = (cmd_channel == 5'b11111);
    assign cmd_is_ts        = (cmd_channel == 5'b10001);
    assign adc_change_mode  = (~prev_cmd_is_ts & cmd_is_ts) | (prev_cmd_is_ts & ~cmd_is_ts);

    always @(posedge clk or negedge rst_n) begin
        if (!rst_n)
            prev_cmd_is_ts  <= 1'b0;
        else if (load_cmd_ready & ~cmd_is_rclb)
            prev_cmd_is_ts  <= cmd_is_ts;
    end

    always @(posedge clk or negedge rst_n) begin
        if (!rst_n)
            cmd_fetched  <= 1'b0;
        else if (load_cmd_fetched)
            cmd_fetched  <= 1'b1;
        else if (clr_cmd_fetched)
            cmd_fetched  <= 1'b0;
    end

    always @(posedge clk or negedge rst_n) begin
        if (!rst_n)
            conv_dly1_s_flp <= 1'b0;
        else
            conv_dly1_s_flp <= conv_dly1_s;
    end

    always @(posedge clk or negedge rst_n) begin
        if (!rst_n)
            pend <= 1'b0;
        else if (conv_dly1_s_flp)
            pend <= 1'b1;
        else if (wait_pend_dly1_s)
            pend <= 1'b0;

    end


    always @(posedge clk or negedge rst_n) begin
        if (!rst_n)
            dout_flp <= 12'd0;
        else if (load_dout)
            dout_flp <= dout;
    end


    always @(posedge clk or negedge rst_n) begin
        if (!rst_n)
            int_timer <= 8'h0;
        else if (load_int_timer)
            int_timer <= 8'h0;
        else if (incr_int_timer)
            int_timer <= int_timer + 8'h1;
    end

    always @(posedge clk or negedge rst_n) begin
        if (!rst_n)
            avrg_cnt_done <= 1'b0;
        else if ((int_timer == (NUM_AVRG_POINTS - 8'd1)) & conv_s)
            avrg_cnt_done <= 1'b1;
        else if (clear_avrg_cnt_done)
            avrg_cnt_done <= 1'b0;
    end

    assign clear_avrg_cnt_done = putresp_dly3_s & ~cmd_valid; // Restart 64 point sampling if continuous sample is broken

    always @(posedge clk or negedge rst_n) begin
        if (!rst_n) begin
            cmd_channel_dly <= 5'h0;
            cmd_sop_dly     <= 1'b0;
            cmd_eop_dly     <= 1'b0;
        end
        else if (load_cmd_ready) begin
            cmd_channel_dly <= cmd_channel;
            cmd_sop_dly     <= cmd_sop;
            cmd_eop_dly     <= cmd_eop;
        end
    end



    assign avrg_enable = cmd_is_ts;

    always @(posedge clk or negedge rst_n) begin
        if (!rst_n)
            avrg_sum    <= 18'h0;
        else if (clear_avrg_sum)
            avrg_sum    <= 18'h0;
        else if (add_avrg_sum_run)
            avrg_sum  <= (avrg_sum - fifo_q) + {6'h0, dout_flp};
        else if (add_avrg_sum)
            avrg_sum  <= avrg_sum + {6'h0, dout_flp};
    end

    assign add_avrg_sum     = ((int_timer != 8'h0) & avrg_cnt_s) |  // when int_timer == 0 the DOUT is not yet ready (ADC hard block introduce one ADC clock delay in the ADC output)
           (conv_dly1_s & avrg_enable & pend) |    // cover averaging pt 64 and beyond (in back 2 back TS scenario)
           (conv_dly1_s & avrg_enable & ~pend & ~frst_64_ptr_done) | // cover averaging pt 63
           (wait_pend_dly1_s & prev_cmd_is_ts); // cover averaging pt 64 and beyond (in switching between ts to non-ts scenario)

    assign add_avrg_sum_run = set_frst_64_ptr_done & frst_64_ptr_done;

    assign clear_avrg_sum           = ~avrg_cnt_done & putresp_pend_s;  // Restart 64 point sampling if continuous sample is broken
    // Not avrg_cnt_done is to ensure put response pending state is caused by broken continuous sampling

    assign set_frst_64_ptr_done     = (wait_pend_dly1_s & prev_cmd_is_ts) | // set at averaging pt 64 and beyond (where next conversion is non-ts)
           (conv_dly1_s & avrg_enable & pend); // set at averaging pt 64 and beyond (where next conversion is ts)
    // No harm to set this signal beyond pt 64

    assign clear_frst_64_ptr_done   = clear_avrg_sum;

    always @(posedge clk or negedge rst_n) begin
        if (!rst_n)
            frst_64_ptr_done <= 1'b0;
        else if (set_frst_64_ptr_done)
            frst_64_ptr_done <= 1'b1;
        else if (clear_frst_64_ptr_done)
            frst_64_ptr_done <= 1'b0;
    end

    assign fifo_sclr    = clear_avrg_sum;
    assign fifo_rdreq   = (((arc_wait_pend_wait_pend_dly1 | arc_sync1_wait_pend_dly1) & prev_cmd_is_ts) | ((arc_conv_conv_dly1 | arc_sync1_conv_dly1) & avrg_enable & pend)) & frst_64_ptr_done;
    assign fifo_wrreq   = ((int_timer != 8'h0) & avrg_cnt_s) |
           (conv_dly1_s & avrg_enable & pend) |
           (conv_dly1_s & avrg_enable & ~pend & ~frst_64_ptr_done) |
           (wait_pend_dly1_s & prev_cmd_is_ts);

    altera_modular_adc_control_avrg_fifo ts_avrg_fifo (
                                             .clock      (clk),
                                             .data       (dout_flp),
                                             .rdreq      (fifo_rdreq),
                                             .wrreq      (fifo_wrreq),
                                             .sclr       (fifo_sclr),
                                             .empty      (),
                                             .full       (),
                                             .q          (fifo_q)
                                         );



    always @(posedge clk or negedge rst_n) begin
        if (!rst_n) begin
            rsp_valid   <= 1'b0;
            rsp_channel <= 5'h0;
            rsp_data    <= 12'h0;
            rsp_sop     <= 1'b0;
            rsp_eop     <= 1'b0;
        end
        else if (load_rsp) begin
            rsp_valid   <= 1'b1;
            rsp_channel <= cmd_channel_dly;
            rsp_data    <= rsp_data_nxt;
            rsp_sop     <= cmd_sop_dly;
            rsp_eop     <= cmd_eop_dly;
        end
        else begin
            rsp_valid   <= 1'b0;
            rsp_channel <= 5'h0;
            rsp_data    <= 12'h0;
            rsp_sop     <= 1'b0;
            rsp_eop     <= 1'b0;
        end
    end

    generate
        if (is_this_first_or_second_adc == 2) begin
            assign rsp_data_nxt = prev_cmd_is_ts ? 12'h0 : dout_flp;    // For ADC2, mask out TSD value since TSD is not supported in ADC2
        end
        else begin
            assign rsp_data_nxt = prev_cmd_is_ts ? avrg_sum[17:6] : dout_flp;
        end
    endgenerate

    always @(posedge clk or negedge rst_n) begin
        if (!rst_n)
            cmd_ready   <= 1'b0;
        else if (load_cmd_ready)
            cmd_ready   <= 1'b1;
        else
            cmd_ready   <= 1'b0;
    end

endmodule




module altera_reset_synchronizer
    #(
         parameter ASYNC_RESET = 1,
         parameter DEPTH       = 2
     )
     (
         input   reset_in /* synthesis ALTERA_ATTRIBUTE = "SUPPRESS_DA_RULE_INTERNAL=R101" */,

         input   clk,
         output  reset_out
     );

    (*preserve*) reg [DEPTH-1:0] altera_reset_synchronizer_int_chain;
    reg altera_reset_synchronizer_int_chain_out;

generate if (ASYNC_RESET) begin
            always @(posedge clk or posedge reset_in) begin
                if (reset_in) begin
                    altera_reset_synchronizer_int_chain <= {DEPTH{1'b1}};
                    altera_reset_synchronizer_int_chain_out <= 1'b1;
                end
                else begin
                    altera_reset_synchronizer_int_chain[DEPTH-2:0] <= altera_reset_synchronizer_int_chain[DEPTH-1:1];
                    altera_reset_synchronizer_int_chain[DEPTH-1] <= 0;
                    altera_reset_synchronizer_int_chain_out <= altera_reset_synchronizer_int_chain[0];
                end
            end

            assign reset_out = altera_reset_synchronizer_int_chain_out;

        end else begin
            always @(posedge clk) begin
                altera_reset_synchronizer_int_chain[DEPTH-2:0] <= altera_reset_synchronizer_int_chain[DEPTH-1:1];
                altera_reset_synchronizer_int_chain[DEPTH-1] <= reset_in;
                altera_reset_synchronizer_int_chain_out <= altera_reset_synchronizer_int_chain[0];
            end

            assign reset_out = altera_reset_synchronizer_int_chain_out;

        end
    endgenerate

endmodule


module fiftyfivenm_adcblock_top_wrapper(
        //reset,               // reset
        chsel,               // 5-bits channel selection.
        soc,                 // signal Start-of-Conversion to ADC
        eoc,                 // signal end of conversion. Data can be latched on the positive edge of clkout_adccore after this signal becomes high.  EOC becomes low at every positive edge of the clkout_adccore signal.
        dout,                // 12-bits DOUT valid after EOC rise, still valid at falling edge, but not before the next EOC rising edge
        usr_pwd,             // User Power Down during run time.  0 = Power Up;  1 = Power Down.
        tsen,                // 0 = Normal Mode; 1 = Temperature Sensing Mode.
        clkout_adccore,      // Output clock from the clock divider
        clkin_from_pll_c0   // Clock source from PLL1 c-counter[0] at BL corner or PLL3 c-counter[0] at TL corner
        //dout_ch              // Indicator to tell that current dout data is for which channel
    );

    // *******************************************************************************************************
    // **   PARAMETERS
    // *******************************************************************************************************

    // -------------------------------------------------------------------------------------------------------
    //      WRAPPED PARAMETERS USED BY fiftyfivenm_adcblock
    // -------------------------------------------------------------------------------------------------------

    // 3-bits 1st stage clock divider.
    // 0..5 = DIV by 1/2/10/20/40/80;
    // 6..7 = invalid
    parameter           clkdiv    = 1;

    // 2nd stage clock divider.
    // 0 = DIV by 10;
    // 1 = DIV by 20
    parameter           tsclkdiv  = 0;

    // 0 = Use 1st stage clock divider when TSEN.
    // 1 = Use 2nd stage clock divider when TSEN.
    parameter           tsclksel  = 0;

    // 2-bits To enable the R ladder for the prescalar input channels.
    // 00 = disable prescalar for CH8 and CH16 (CH8 for device with 2nd ADC)
    // 01 = enable prescalar for CH8 only
    // 10 = enable prescalar for CH16 only (CH8 for device with 2nd ADC)
    // 11 = enable prescalar for CH8 and CH16 (CH8 for device with 2nd ADC)
    // please note that this is not supported in VR mode
    parameter           prescalar = 0;

    // Reference voltage selection for ADC.
    // 0 = external;
    // 1 = internal VCCADC_2P5
    parameter           refsel    = 0;

    // -------------------------------------------------------------------------------------------------------
    //      WRAPPED PARAMETERS  USED BY both chsel_code_converter_sw_to_hw and fiftyfivenm_adcblock
    // -------------------------------------------------------------------------------------------------------

    // Ordering Part Number 10MXX... code
    parameter           device_partname_fivechar_prefix = "10M08";      // Valid options = 04, 08, 16, 25, 40, 50

    // Some part have two ADC, instantiate which ADC?  1st or 2nd?
    parameter           is_this_first_or_second_adc = 1;    // Valid options = 1 or 2

    // 16 bits to indicate whether each of the dual purpose analog input pin (ADCIN) is in use or not.
    // 1 bit to indicate whether dedicated analog input pin (ANAIN) is in use or not (bit 16)
    parameter           analog_input_pin_mask = 17'h0;

    // Power Down. Use to disable the ADC during compilation time if no ADC is in use.
    parameter           hard_pwd = 0;

    // Logic simulation parameters which only affects simulation behavior
    parameter           enable_usr_sim = 0;
    parameter           reference_voltage_sim = 65536;
    parameter           simfilename_ch0 = "simfilename_ch0";
    parameter           simfilename_ch1 = "simfilename_ch1";
    parameter           simfilename_ch2 = "simfilename_ch2";
    parameter           simfilename_ch3 = "simfilename_ch3";
    parameter           simfilename_ch4 = "simfilename_ch4";
    parameter           simfilename_ch5 = "simfilename_ch5";
    parameter           simfilename_ch6 = "simfilename_ch6";
    parameter           simfilename_ch7 = "simfilename_ch7";
    parameter           simfilename_ch8 = "simfilename_ch8";
    parameter           simfilename_ch9 = "simfilename_ch9";
    parameter           simfilename_ch10 = "simfilename_ch10";
    parameter           simfilename_ch11 = "simfilename_ch11";
    parameter           simfilename_ch12 = "simfilename_ch12";
    parameter           simfilename_ch13 = "simfilename_ch13";
    parameter           simfilename_ch14 = "simfilename_ch14";
    parameter           simfilename_ch15 = "simfilename_ch15";
    parameter           simfilename_ch16 = "simfilename_ch16";

    // *******************************************************************************************************
    // **   INPUTS
    // *******************************************************************************************************

    //input               reset;      // reset

    input               clkin_from_pll_c0;  // Clock source from PLL1 c-counter[0] at BL corner or PLL3 c-counter[0] at TL corner

    input               soc;        // signal Start-of-Conversion to ADC
    input               usr_pwd;    // User Power Down during run time.  0 = Power Up;  1 = Power Down.
    input               tsen;       // 0 = Normal Mode; 1 = Temperature Sensing Mode.
    input   [4:0]       chsel;      // 5-bits channel selection.

    // *******************************************************************************************************
    // **   OUTPUTS
    // *******************************************************************************************************

    output              clkout_adccore;  // Output clock from the clock divider
    output              eoc;        // signal end of conversion. Data can be latched on the positive edge of clkout_adccore after this signal becomes high.  EOC becomes low at every positive edge of the clkout_adccore signal.
    output [11:0]       dout;       // 12-bits DOUT valid after EOC rise, still valid at falling edge, but not before the next EOC rising edge
    wire    [4:0]       chsel_to_hw;

    chsel_code_converter_sw_to_hw decoder(
                                      // The 5-bits chsel input port are wired to chsel_from_sw for conversion
                                      .chsel_from_sw(chsel),
                                      // The chsel_code_converter_sw_to_hw output chsel_to_hw which will be wired into fiftyfivenm_adcblock
                                      .chsel_to_hw(chsel_to_hw)
                                  );
    defparam           decoder.device_partname_fivechar_prefix = device_partname_fivechar_prefix;
    defparam           decoder.is_this_first_or_second_adc     = is_this_first_or_second_adc;

    // -------------------------------------------------------------------------------------------------------
    //      2.00: Instantiate ADC Block primitive
    // -------------------------------------------------------------------------------------------------------

    fiftyfivenm_adcblock_primitive_wrapper adcblock_instance(
                                               // .reset            (reset),
                                               .chsel            (chsel_to_hw),
                                               .soc              (soc),
                                               .eoc              (eoc),
                                               .dout             (dout),
                                               .usr_pwd          (usr_pwd),
                                               .tsen             (tsen),
                                               .clkout_adccore   (clkout_adccore),
                                               .clkin_from_pll_c0(clkin_from_pll_c0)
                                           );
    defparam  adcblock_instance.clkdiv                          = clkdiv;
    defparam  adcblock_instance.tsclkdiv                        = tsclkdiv;
    defparam  adcblock_instance.tsclksel                        = tsclksel;
    defparam  adcblock_instance.prescalar                       = prescalar;
    defparam  adcblock_instance.refsel                          = refsel;
    defparam  adcblock_instance.device_partname_fivechar_prefix = device_partname_fivechar_prefix;
    defparam  adcblock_instance.is_this_first_or_second_adc     = is_this_first_or_second_adc;
    defparam  adcblock_instance.analog_input_pin_mask           = analog_input_pin_mask;
    defparam  adcblock_instance.hard_pwd                        = hard_pwd;
    defparam  adcblock_instance.enable_usr_sim                  = enable_usr_sim;
    defparam  adcblock_instance.reference_voltage_sim           = reference_voltage_sim;
    defparam  adcblock_instance.simfilename_ch0                 = simfilename_ch0;
    defparam  adcblock_instance.simfilename_ch1                 = simfilename_ch1;
    defparam  adcblock_instance.simfilename_ch2                 = simfilename_ch2;
    defparam  adcblock_instance.simfilename_ch3                 = simfilename_ch3;
    defparam  adcblock_instance.simfilename_ch4                 = simfilename_ch4;
    defparam  adcblock_instance.simfilename_ch5                 = simfilename_ch5;
    defparam  adcblock_instance.simfilename_ch6                 = simfilename_ch6;
    defparam  adcblock_instance.simfilename_ch7                 = simfilename_ch7;
    defparam  adcblock_instance.simfilename_ch8                 = simfilename_ch8;
    defparam  adcblock_instance.simfilename_ch9                 = simfilename_ch9;
    defparam  adcblock_instance.simfilename_ch10                = simfilename_ch10;
    defparam  adcblock_instance.simfilename_ch11                = simfilename_ch11;
    defparam  adcblock_instance.simfilename_ch12                = simfilename_ch12;
    defparam  adcblock_instance.simfilename_ch13                = simfilename_ch13;
    defparam  adcblock_instance.simfilename_ch14                = simfilename_ch14;
    defparam  adcblock_instance.simfilename_ch15                = simfilename_ch15;
    defparam  adcblock_instance.simfilename_ch16                = simfilename_ch16;

endmodule

module altera_reset_controller
    #(
         parameter NUM_RESET_INPUTS              = 6,
         parameter USE_RESET_REQUEST_IN0 = 0,
         parameter USE_RESET_REQUEST_IN1 = 0,
         parameter USE_RESET_REQUEST_IN2 = 0,
         parameter USE_RESET_REQUEST_IN3 = 0,
         parameter USE_RESET_REQUEST_IN4 = 0,
         parameter USE_RESET_REQUEST_IN5 = 0,
         parameter USE_RESET_REQUEST_IN6 = 0,
         parameter USE_RESET_REQUEST_IN7 = 0,
         parameter USE_RESET_REQUEST_IN8 = 0,
         parameter USE_RESET_REQUEST_IN9 = 0,
         parameter USE_RESET_REQUEST_IN10 = 0,
         parameter USE_RESET_REQUEST_IN11 = 0,
         parameter USE_RESET_REQUEST_IN12 = 0,
         parameter USE_RESET_REQUEST_IN13 = 0,
         parameter USE_RESET_REQUEST_IN14 = 0,
         parameter USE_RESET_REQUEST_IN15 = 0,
         parameter OUTPUT_RESET_SYNC_EDGES       = "deassert",
         parameter SYNC_DEPTH                    = 2,
         parameter RESET_REQUEST_PRESENT         = 0,
         parameter RESET_REQ_WAIT_TIME           = 3,
         parameter MIN_RST_ASSERTION_TIME        = 11,
         parameter RESET_REQ_EARLY_DSRT_TIME     = 4,
         parameter ADAPT_RESET_REQUEST          = 0
     )
     (
         // --------------------------------------
         // We support up to 16 reset inputs, for now
         // --------------------------------------
         input reset_in0,
         input reset_in1,
         input reset_in2,
         input reset_in3,
         input reset_in4,
         input reset_in5,
         input reset_in6,
         input reset_in7,
         input reset_in8,
         input reset_in9,
         input reset_in10,
         input reset_in11,
         input reset_in12,
         input reset_in13,
         input reset_in14,
         input reset_in15,
         input reset_req_in0,
         input reset_req_in1,
         input reset_req_in2,
         input reset_req_in3,
         input reset_req_in4,
         input reset_req_in5,
         input reset_req_in6,
         input reset_req_in7,
         input reset_req_in8,
         input reset_req_in9,
         input reset_req_in10,
         input reset_req_in11,
         input reset_req_in12,
         input reset_req_in13,
         input reset_req_in14,
         input reset_req_in15,


         input  clk,
         output reg reset_out,
         output reg reset_req
     );

    // Always use async reset synchronizer if reset_req is used
    localparam ASYNC_RESET = (OUTPUT_RESET_SYNC_EDGES == "deassert");

    // --------------------------------------
    // Local parameter to control the reset_req and reset_out timing when RESET_REQUEST_PRESENT==1
    // --------------------------------------
    localparam MIN_METASTABLE = 3;
    localparam RSTREQ_ASRT_SYNC_TAP = MIN_METASTABLE + RESET_REQ_WAIT_TIME;

    localparam LARGER = RESET_REQ_WAIT_TIME > RESET_REQ_EARLY_DSRT_TIME ? RESET_REQ_WAIT_TIME : RESET_REQ_EARLY_DSRT_TIME;

    localparam ASSERTION_CHAIN_LENGTH =  (MIN_METASTABLE > LARGER) ?
               MIN_RST_ASSERTION_TIME + 1 :
               (
                   (MIN_RST_ASSERTION_TIME > LARGER)?
                   MIN_RST_ASSERTION_TIME + (LARGER - MIN_METASTABLE + 1) + 1 :
                   MIN_RST_ASSERTION_TIME + RESET_REQ_EARLY_DSRT_TIME + RESET_REQ_WAIT_TIME - MIN_METASTABLE + 2
               );

    localparam RESET_REQ_DRST_TAP = RESET_REQ_EARLY_DSRT_TIME + 1;
    // --------------------------------------

    wire merged_reset;
    wire merged_reset_req_in;
    wire reset_out_pre;
    wire reset_req_pre;

    // Registers and Interconnect
    (*preserve*) reg  [RSTREQ_ASRT_SYNC_TAP: 0]  altera_reset_synchronizer_int_chain;
    reg [ASSERTION_CHAIN_LENGTH-1: 0]            r_sync_rst_chain;
    reg                                          r_sync_rst;
    reg                                          r_early_rst;

    // --------------------------------------
    // "Or" all the input resets together
    // --------------------------------------
    assign merged_reset = (
               reset_in0 |
               reset_in1 |
               reset_in2 |
               reset_in3 |
               reset_in4 |
               reset_in5 |
               reset_in6 |
               reset_in7 |
               reset_in8 |
               reset_in9 |
               reset_in10 |
               reset_in11 |
               reset_in12 |
               reset_in13 |
               reset_in14 |
               reset_in15
           );

    assign merged_reset_req_in = (
               ( (USE_RESET_REQUEST_IN0 == 1) ? reset_req_in0 : 1'b0)  |
               ( (USE_RESET_REQUEST_IN1 == 1) ? reset_req_in1 : 1'b0)  |
               ( (USE_RESET_REQUEST_IN2 == 1) ? reset_req_in2 : 1'b0)  |
               ( (USE_RESET_REQUEST_IN3 == 1) ? reset_req_in3 : 1'b0)  |
               ( (USE_RESET_REQUEST_IN4 == 1) ? reset_req_in4 : 1'b0)  |
               ( (USE_RESET_REQUEST_IN5 == 1) ? reset_req_in5 : 1'b0)  |
               ( (USE_RESET_REQUEST_IN6 == 1) ? reset_req_in6 : 1'b0)  |
               ( (USE_RESET_REQUEST_IN7 == 1) ? reset_req_in7 : 1'b0)  |
               ( (USE_RESET_REQUEST_IN8 == 1) ? reset_req_in8 : 1'b0)  |
               ( (USE_RESET_REQUEST_IN9 == 1) ? reset_req_in9 : 1'b0)  |
               ( (USE_RESET_REQUEST_IN10 == 1) ? reset_req_in10 : 1'b0)  |
               ( (USE_RESET_REQUEST_IN11 == 1) ? reset_req_in11 : 1'b0)  |
               ( (USE_RESET_REQUEST_IN12 == 1) ? reset_req_in12 : 1'b0)  |
               ( (USE_RESET_REQUEST_IN13 == 1) ? reset_req_in13 : 1'b0)  |
               ( (USE_RESET_REQUEST_IN14 == 1) ? reset_req_in14 : 1'b0)  |
               ( (USE_RESET_REQUEST_IN15 == 1) ? reset_req_in15 : 1'b0)
           );


    // --------------------------------------
    // And if required, synchronize it to the required clock domain,
    // with the correct synchronization type
    // --------------------------------------
generate if (OUTPUT_RESET_SYNC_EDGES == "none" && (RESET_REQUEST_PRESENT==0)) begin

            assign reset_out_pre = merged_reset;
            assign reset_req_pre = merged_reset_req_in;

        end else begin

            altera_reset_synchronizer
                #(
                    .DEPTH      (SYNC_DEPTH),
                    .ASYNC_RESET(RESET_REQUEST_PRESENT? 1'b1 : ASYNC_RESET)
                )
                alt_rst_sync_uq1
                (
                    .clk        (clk),
                    .reset_in   (merged_reset),
                    .reset_out  (reset_out_pre)
                );

            altera_reset_synchronizer
                #(
                    .DEPTH      (SYNC_DEPTH),
                    .ASYNC_RESET(0)
                )
                alt_rst_req_sync_uq1
                (
                    .clk        (clk),
                    .reset_in   (merged_reset_req_in),
                    .reset_out  (reset_req_pre)
                );

        end
    endgenerate

    generate if ( ( (RESET_REQUEST_PRESENT == 0) && (ADAPT_RESET_REQUEST==0) )|
                      ( (ADAPT_RESET_REQUEST == 1) && (OUTPUT_RESET_SYNC_EDGES != "deassert") ) ) begin
            always @* begin
                reset_out = reset_out_pre;
                reset_req = reset_req_pre;
            end
        end else if ( (RESET_REQUEST_PRESENT == 0) && (ADAPT_RESET_REQUEST==1) ) begin

            wire reset_out_pre2;

            altera_reset_synchronizer
                #(
                    .DEPTH      (SYNC_DEPTH+1),
                    .ASYNC_RESET(0)
                )
                alt_rst_sync_uq2
                (
                    .clk        (clk),
                    .reset_in   (reset_out_pre),
                    .reset_out  (reset_out_pre2)
                );

            always @* begin
                reset_out = reset_out_pre2;
                reset_req = reset_req_pre;
            end

        end
        else begin

            // 3-FF Metastability Synchronizer
            initial
            begin
                altera_reset_synchronizer_int_chain <= {RSTREQ_ASRT_SYNC_TAP{1'b1}};
            end

            always @(posedge clk)
            begin
                altera_reset_synchronizer_int_chain[RSTREQ_ASRT_SYNC_TAP:0] <=
                                                   {altera_reset_synchronizer_int_chain[RSTREQ_ASRT_SYNC_TAP-1:0], reset_out_pre};
            end

            // Synchronous reset pipe
            initial
            begin
                r_sync_rst_chain <= {ASSERTION_CHAIN_LENGTH{1'b1}};
            end

            always @(posedge clk)
            begin
                if (altera_reset_synchronizer_int_chain[MIN_METASTABLE-1] == 1'b1)
                begin
                    r_sync_rst_chain <= {ASSERTION_CHAIN_LENGTH{1'b1}};
                end
                else
                begin
                    r_sync_rst_chain <= {1'b0, r_sync_rst_chain[ASSERTION_CHAIN_LENGTH-1:1]};
                end
            end

            // Standard synchronous reset output.  From 0-1, the transition lags the early output.  For 1->0, the transition
            // matches the early input.

            always @(posedge clk)
            begin
                case ({altera_reset_synchronizer_int_chain[RSTREQ_ASRT_SYNC_TAP], r_sync_rst_chain[1], r_sync_rst})
                    3'b000:   r_sync_rst <= 1'b0; // Not reset
                    3'b001:   r_sync_rst <= 1'b0;
                    3'b010:   r_sync_rst <= 1'b0;
                    3'b011:   r_sync_rst <= 1'b1;
                    3'b100:   r_sync_rst <= 1'b1;
                    3'b101:   r_sync_rst <= 1'b1;
                    3'b110:   r_sync_rst <= 1'b1;
                    3'b111:   r_sync_rst <= 1'b1; // In Reset
                    default:  r_sync_rst <= 1'b1;
                endcase

                case ({r_sync_rst_chain[1], r_sync_rst_chain[RESET_REQ_DRST_TAP] | reset_req_pre})
                    2'b00:   r_early_rst <= 1'b0; // Not reset
                    2'b01:   r_early_rst <= 1'b1; // Coming out of reset
                    2'b10:   r_early_rst <= 1'b0; // Spurious reset - should not be possible via synchronous design.
                    2'b11:   r_early_rst <= 1'b1; // Held in reset
                    default: r_early_rst <= 1'b1;
                endcase
            end

            always @* begin
                reset_out = r_sync_rst;
                reset_req = r_early_rst;
            end

        end
    endgenerate

endmodule




module altera_modular_adc_control_avrg_fifo (
        clock,
        data,
        rdreq,
        sclr,
        wrreq,
        empty,
        full,
        q);

    input	  clock;
    input	[11:0]  data;
    input	  rdreq;
    input	  sclr;
    input	  wrreq;
    output	  empty;
    output	  full;
    output	[11:0]  q;

    wire  sub_wire0;
    wire  sub_wire1;
    wire [11:0] sub_wire2;
    wire  empty = sub_wire0;
    wire  full = sub_wire1;
    wire [11:0] q = sub_wire2[11:0];

    scfifo	scfifo_component (
               .clock (clock),
               .data (data),
               .rdreq (rdreq),
               .sclr (sclr),
               .wrreq (wrreq),
               .empty (sub_wire0),
               .full (sub_wire1),
               .q (sub_wire2),
               .aclr (),
               .almost_empty (),
               .almost_full (),
               .usedw ());
    defparam
        scfifo_component.add_ram_output_register = "OFF",
        scfifo_component.intended_device_family = "MAX 10",
        scfifo_component.lpm_hint = "RAM_BLOCK_TYPE=M9K",
        scfifo_component.lpm_numwords = 64,
        scfifo_component.lpm_showahead = "OFF",
        scfifo_component.lpm_type = "scfifo",
        scfifo_component.lpm_width = 12,
        scfifo_component.lpm_widthu = 6,
        scfifo_component.overflow_checking = "ON",
        scfifo_component.underflow_checking = "ON",
        scfifo_component.use_eab = "ON";

endmodule


module  chsel_code_converter_sw_to_hw (
        chsel_from_sw,            // 5-bits channel selection.
        chsel_to_hw               // 5-bits channel selection.
    );

    parameter           device_partname_fivechar_prefix = "10M08";   // Valid options = 04, 08, 16, 25, 40, 50
    parameter           is_this_first_or_second_adc = 1;             // Valid options = 1 or 2
    localparam          variant_08n16_hw_chsel_code_for_sw_temp_code_10001 = 5'b00000;
    localparam          variant_08n16_hw_chsel_code_for_sw_ch00_code_00000 = 5'b00011;
    localparam          variant_08n16_hw_chsel_code_for_sw_ch01_code_00001 = 5'b00100;
    localparam          variant_08n16_hw_chsel_code_for_sw_ch02_code_00010 = 5'b00110;
    localparam          variant_08n16_hw_chsel_code_for_sw_ch03_code_00011 = 5'b01010;
    localparam          variant_08n16_hw_chsel_code_for_sw_ch04_code_00100 = 5'b01100;
    localparam          variant_08n16_hw_chsel_code_for_sw_ch05_code_00101 = 5'b10000;
    localparam          variant_08n16_hw_chsel_code_for_sw_ch06_code_00110 = 5'b01110;
    localparam          variant_08n16_hw_chsel_code_for_sw_ch07_code_00111 = 5'b01101;
    localparam          variant_08n16_hw_chsel_code_for_sw_ch08_code_01000 = 5'b00010;
    localparam          variant_08n16_hw_chsel_code_for_sw_ch09_code_01001 = 5'b00101;
    localparam          variant_08n16_hw_chsel_code_for_sw_ch10_code_01010 = 5'b01001;
    localparam          variant_08n16_hw_chsel_code_for_sw_ch11_code_01011 = 5'b10001;
    localparam          variant_08n16_hw_chsel_code_for_sw_ch12_code_01100 = 5'b01111;
    localparam          variant_08n16_hw_chsel_code_for_sw_ch13_code_01101 = 5'b01000;
    localparam          variant_08n16_hw_chsel_code_for_sw_ch14_code_01110 = 5'b00111;
    localparam          variant_08n16_hw_chsel_code_for_sw_ch15_code_01111 = 5'b01011;
    localparam          variant_08n16_hw_chsel_code_for_sw_ch16_code_10000 = 5'b00001;

    // First ADC of 10M25/40/50 hardware equivalent chsel code for a particular software chsel code
    localparam          dual_first_adc_hw_chsel_code_for_sw_temp_code_10001 = 5'b00000;
    localparam          dual_first_adc_hw_chsel_code_for_sw_ch00_code_00000 = 5'b00011;
    localparam          dual_first_adc_hw_chsel_code_for_sw_ch01_code_00001 = 5'b00100;
    localparam          dual_first_adc_hw_chsel_code_for_sw_ch02_code_00010 = 5'b00110;
    localparam          dual_first_adc_hw_chsel_code_for_sw_ch03_code_00011 = 5'b01010;
    localparam          dual_first_adc_hw_chsel_code_for_sw_ch04_code_00100 = 5'b01100;
    localparam          dual_first_adc_hw_chsel_code_for_sw_ch05_code_00101 = 5'b10000;
    localparam          dual_first_adc_hw_chsel_code_for_sw_ch06_code_00110 = 5'b01110;
    localparam          dual_first_adc_hw_chsel_code_for_sw_ch07_code_00111 = 5'b01101;
    localparam          dual_first_adc_hw_chsel_code_for_sw_ch08_code_01000 = 5'b00010;

    // Second ADC of 10M25/40/50 hardware equivalent chsel code for a particular software chsel code
    // Note that: Second ADC do not support internal temperature sensor.
    // However internal temperature sensor mapping for ADC2 is later included for dual adc mode
    // When in dual adc mode, if ADC1 is operating in TSD mode, ADC2 will perform a dummy TSD mode as well
    localparam          dual_second_adc_hw_chsel_code_for_sw_temp_code_10001 = 5'b00000;
    localparam          dual_second_adc_hw_chsel_code_for_sw_ch00_code_00000 = 5'b00011;
    localparam          dual_second_adc_hw_chsel_code_for_sw_ch01_code_00001 = 5'b00101;
    localparam          dual_second_adc_hw_chsel_code_for_sw_ch02_code_00010 = 5'b01001;
    localparam          dual_second_adc_hw_chsel_code_for_sw_ch03_code_00011 = 5'b10001;
    localparam          dual_second_adc_hw_chsel_code_for_sw_ch04_code_00100 = 5'b01111;
    localparam          dual_second_adc_hw_chsel_code_for_sw_ch05_code_00101 = 5'b01000;
    localparam          dual_second_adc_hw_chsel_code_for_sw_ch06_code_00110 = 5'b00111;
    localparam          dual_second_adc_hw_chsel_code_for_sw_ch07_code_00111 = 5'b01011;
    localparam          dual_second_adc_hw_chsel_code_for_sw_ch08_code_01000 = 5'b00001;

    // *******************************************************************************************************
    // **   INPUTS
    // *******************************************************************************************************

    input   [4:0]       chsel_from_sw;  // 5-bits channel selection number from software perspective

    // *******************************************************************************************************
    // **   OUTPUTS
    // *******************************************************************************************************

    output  [4:0]       chsel_to_hw;    // 5-bits channel selection code to be send to ADC Hard IP

    // *******************************************************************************************************
    // **   EXTERNAL NET AND REGISTER DATA TYPE (with input / output / inout ports)
    // *******************************************************************************************************

    reg     [4:0]       chsel_to_hw;    // 5-bits channel selection code to be send to ADC Hard IP

    // *******************************************************************************************************
    // **   MAIN CODE
    // *******************************************************************************************************

    // -------------------------------------------------------------------------------------------------------
    //      1.00: Channel Mapping
    // -------------------------------------------------------------------------------------------------------

    // DESCRIBE THE ALWAYS BLOCK:
    // This block execute on divided internal clock
    // Its job is mainly to determine what value to be set for the digital_out and eoc_rise
    always @(chsel_from_sw)
    begin
        // DESCRIBE THE CASE STATEMENT:
        // Output the equivalent chsel code for hardware
        if  ((device_partname_fivechar_prefix == "10M04") || (device_partname_fivechar_prefix == "10M08") || (device_partname_fivechar_prefix == "10M16"))
        begin
            // COMMENT FOR THIS BRANCH:
            // 10M08/04 channel mapping
            case(chsel_from_sw)
                5'b10001: chsel_to_hw <= variant_08n16_hw_chsel_code_for_sw_temp_code_10001;
                5'b00000: chsel_to_hw <= variant_08n16_hw_chsel_code_for_sw_ch00_code_00000;
                5'b00001: chsel_to_hw <= variant_08n16_hw_chsel_code_for_sw_ch01_code_00001;
                5'b00010: chsel_to_hw <= variant_08n16_hw_chsel_code_for_sw_ch02_code_00010;
                5'b00011: chsel_to_hw <= variant_08n16_hw_chsel_code_for_sw_ch03_code_00011;
                5'b00100: chsel_to_hw <= variant_08n16_hw_chsel_code_for_sw_ch04_code_00100;
                5'b00101: chsel_to_hw <= variant_08n16_hw_chsel_code_for_sw_ch05_code_00101;
                5'b00110: chsel_to_hw <= variant_08n16_hw_chsel_code_for_sw_ch06_code_00110;
                5'b00111: chsel_to_hw <= variant_08n16_hw_chsel_code_for_sw_ch07_code_00111;
                5'b01000: chsel_to_hw <= variant_08n16_hw_chsel_code_for_sw_ch08_code_01000;
                5'b01001: chsel_to_hw <= variant_08n16_hw_chsel_code_for_sw_ch09_code_01001;
                5'b01010: chsel_to_hw <= variant_08n16_hw_chsel_code_for_sw_ch10_code_01010;
                5'b01011: chsel_to_hw <= variant_08n16_hw_chsel_code_for_sw_ch11_code_01011;
                5'b01100: chsel_to_hw <= variant_08n16_hw_chsel_code_for_sw_ch12_code_01100;
                5'b01101: chsel_to_hw <= variant_08n16_hw_chsel_code_for_sw_ch13_code_01101;
                5'b01110: chsel_to_hw <= variant_08n16_hw_chsel_code_for_sw_ch14_code_01110;
                5'b01111: chsel_to_hw <= variant_08n16_hw_chsel_code_for_sw_ch15_code_01111;
                5'b10000: chsel_to_hw <= variant_08n16_hw_chsel_code_for_sw_ch16_code_10000;
                default : chsel_to_hw <= 5'b11111;
            endcase
        end
        else
            if ((is_this_first_or_second_adc == 1) &&
                    ((device_partname_fivechar_prefix == "10M25") ||
                     (device_partname_fivechar_prefix == "10M40") ||
                     (device_partname_fivechar_prefix == "10M50")))
            begin
                // COMMENT FOR THIS BRANCH:
                // First ADC of 10M25/40/50 channel mapping
                case(chsel_from_sw)
                    5'b10001: chsel_to_hw <= dual_first_adc_hw_chsel_code_for_sw_temp_code_10001;
                    5'b00000: chsel_to_hw <= dual_first_adc_hw_chsel_code_for_sw_ch00_code_00000;
                    5'b00001: chsel_to_hw <= dual_first_adc_hw_chsel_code_for_sw_ch01_code_00001;
                    5'b00010: chsel_to_hw <= dual_first_adc_hw_chsel_code_for_sw_ch02_code_00010;
                    5'b00011: chsel_to_hw <= dual_first_adc_hw_chsel_code_for_sw_ch03_code_00011;
                    5'b00100: chsel_to_hw <= dual_first_adc_hw_chsel_code_for_sw_ch04_code_00100;
                    5'b00101: chsel_to_hw <= dual_first_adc_hw_chsel_code_for_sw_ch05_code_00101;
                    5'b00110: chsel_to_hw <= dual_first_adc_hw_chsel_code_for_sw_ch06_code_00110;
                    5'b00111: chsel_to_hw <= dual_first_adc_hw_chsel_code_for_sw_ch07_code_00111;
                    5'b01000: chsel_to_hw <= dual_first_adc_hw_chsel_code_for_sw_ch08_code_01000;
                    default : chsel_to_hw <= 5'b11111;
                endcase
            end
            else
                if ((is_this_first_or_second_adc == 2) &&
                        ((device_partname_fivechar_prefix == "10M25") ||
                         (device_partname_fivechar_prefix == "10M40") ||
                         (device_partname_fivechar_prefix == "10M50")))
                begin
                    // COMMENT FOR THIS BRANCH:
                    // Second ADC of 10M25/40/50 channel mapping
                    case(chsel_from_sw)
                        5'b10001: chsel_to_hw <= dual_second_adc_hw_chsel_code_for_sw_temp_code_10001;
                        5'b00000: chsel_to_hw <= dual_second_adc_hw_chsel_code_for_sw_ch00_code_00000;
                        5'b00001: chsel_to_hw <= dual_second_adc_hw_chsel_code_for_sw_ch01_code_00001;
                        5'b00010: chsel_to_hw <= dual_second_adc_hw_chsel_code_for_sw_ch02_code_00010;
                        5'b00011: chsel_to_hw <= dual_second_adc_hw_chsel_code_for_sw_ch03_code_00011;
                        5'b00100: chsel_to_hw <= dual_second_adc_hw_chsel_code_for_sw_ch04_code_00100;
                        5'b00101: chsel_to_hw <= dual_second_adc_hw_chsel_code_for_sw_ch05_code_00101;
                        5'b00110: chsel_to_hw <= dual_second_adc_hw_chsel_code_for_sw_ch06_code_00110;
                        5'b00111: chsel_to_hw <= dual_second_adc_hw_chsel_code_for_sw_ch07_code_00111;
                        5'b01000: chsel_to_hw <= dual_second_adc_hw_chsel_code_for_sw_ch08_code_01000;
                        default : chsel_to_hw <= 5'b11111;
                    endcase
                end
    end // end always

endmodule



module fiftyfivenm_adcblock_primitive_wrapper(
        //reset,
        chsel,               // 5-bits channel selection.
        soc,                 // signal Start-of-Conversion to ADC
        eoc,                 // signal end of conversion. Data can be latched on the positive edge of clk_dft after this signal becomes high.  EOC becomes low at every positive edge of the clk_dft signal.
        dout,                // 12-bits DOUT valid after EOC rise, still valid at falling edge, but not before the next EOC rising edge
        usr_pwd,             // User Power Down during run time.  0 = Power Up;  1 = Power Down.
        tsen,                // 0 = Normal Mode; 1 = Temperature Sensing Mode.
        clkout_adccore,      // Output clock from the clock divider
        clkin_from_pll_c0    // Clock source from PLL1 c-counter[0] at BL corner or PLL3 c-counter[0] at TL corner
    );

    // *******************************************************************************************************
    // **   PARAMETERS
    // *******************************************************************************************************

    // -------------------------------------------------------------------------------------------------------
    //      WRAPPED PARAMETERS USED BY fiftyfivenm_adcblock
    // -------------------------------------------------------------------------------------------------------

    // 3-bits 1st stage clock divider.
    // 0..5 = DIV by 1/2/10/20/40/80;
    // 6..7 = invalid
    parameter           clkdiv    = 1;

    // 2nd stage clock divider.
    // 0 = DIV by 10;
    // 1 = DIV by 20
    parameter           tsclkdiv  = 0;

    // 0 = Use 1st stage clock divider when TSEN.
    // 1 = Use 2nd stage clock divider when TSEN.
    parameter           tsclksel  = 0;

    // 2-bits To enable the R ladder for the prescalar input channels.
    // 00 = disable prescalar for CH8 and CH16 (CH8 for device with 2nd ADC)
    // 01 = enable prescalar for CH8 only
    // 10 = enable prescalar for CH16 only (CH8 for device with 2nd ADC)
    // 11 = enable prescalar for CH8 and CH16 (CH8 for device with 2nd ADC)
    // please note that this is not supported in VR mode
    parameter           prescalar = 0;

    // Reference voltage selection for ADC.
    // 0 = external;
    // 1 = internal VCCADC_2P5
    parameter           refsel    = 0;

    // Ordering Part Number 10MXX... code
    parameter           device_partname_fivechar_prefix = "10M08";      // Valid options = 04, 08, 16, 25, 40, 50

    // Some part have two ADC, instantiate which ADC?  1st or 2nd?
    parameter           is_this_first_or_second_adc = 1;    // Valid options = 1 or 2

    // is_using_dedicated_analog_input_pin_only? -> removed, replaced with analog_input_pin_mask
    //parameter           is_using_dedicated_analog_input_pin_only = 0;

    // 16 bits to indicate whether each of the dual purpose analog input pin (ADCIN) is in use or not.
    // 1 bit to indicate whether dedicated analog input pin (ANAIN) is in use or not (bit 16)
    parameter           analog_input_pin_mask = 17'h0;

    // Power Down. Use to disable the ADC during compilation time if no ADC is in use.
    parameter           hard_pwd = 0;

    // Logic simulation parameters which only affects simulation behavior
    parameter           enable_usr_sim = 0;
    parameter           reference_voltage_sim = 65536;
    parameter           simfilename_ch0 = "simfilename_ch0";
    parameter           simfilename_ch1 = "simfilename_ch1";
    parameter           simfilename_ch2 = "simfilename_ch2";
    parameter           simfilename_ch3 = "simfilename_ch3";
    parameter           simfilename_ch4 = "simfilename_ch4";
    parameter           simfilename_ch5 = "simfilename_ch5";
    parameter           simfilename_ch6 = "simfilename_ch6";
    parameter           simfilename_ch7 = "simfilename_ch7";
    parameter           simfilename_ch8 = "simfilename_ch8";
    parameter           simfilename_ch9 = "simfilename_ch9";
    parameter           simfilename_ch10 = "simfilename_ch10";
    parameter           simfilename_ch11 = "simfilename_ch11";
    parameter           simfilename_ch12 = "simfilename_ch12";
    parameter           simfilename_ch13 = "simfilename_ch13";
    parameter           simfilename_ch14 = "simfilename_ch14";
    parameter           simfilename_ch15 = "simfilename_ch15";
    parameter           simfilename_ch16 = "simfilename_ch16";


    // *******************************************************************************************************
    // **   INPUTS
    // *******************************************************************************************************

    //input               reset;

    input               clkin_from_pll_c0;  // Clock source from PLL1 c-counter[0] at BL corner or PLL3 c-counter[0] at TL corner

    input               soc;        // signal Start-of-Conversion to ADC
    input               usr_pwd;    // User Power Down during run time.  0 = Power Up;  1 = Power Down.
    input               tsen;       // 0 = Normal Mode; 1 = Temperature Sensing Mode.
    input   [4:0]       chsel;      // 5-bits channel selection.

    //reg                 reg_clk_dft_soc;
    //reg     [4:0]       reg_clk_dft_chsel;

    // *******************************************************************************************************
    // **   OUTPUTS
    // *******************************************************************************************************

    output              clkout_adccore;
    output              eoc;

    output  [11:0]      dout;
    wire    [11:0]      wire_from_adc_dout;
    //reg     [11:0]      reg_clk_dft_dout;

    // *******************************************************************************************************
    // **   OUTPUTS ASSIGNMENTS
    // *******************************************************************************************************

    //assign       dout = reg_clk_dft_dout;
    assign       dout = wire_from_adc_dout;

    // *******************************************************************************************************
    // **   INITIALIZATION
    // *******************************************************************************************************

    // *******************************************************************************************************
    // **   MAIN CODE
    // *******************************************************************************************************

    // -------------------------------------------------------------------------------------------------------
    //      1.00: Instantiate ADC Block primitive
    // -------------------------------------------------------------------------------------------------------
`ifdef DEBUG_AND_DEVELOPMENT
    fiftyfivenm_adcblock_emulation primitive_instance(
`else
    fiftyfivenm_adcblock primitive_instance(
`endif
                                       //.chsel            (reg_clk_dft_chsel),
                                       //.soc              (reg_clk_dft_soc),
                                       .chsel            (chsel),
                                       .soc              (soc),
                                       .eoc              (eoc),
                                       .dout             (wire_from_adc_dout),
                                       .usr_pwd          (usr_pwd),
                                       .tsen             (tsen),
                                       .clk_dft          (clkout_adccore),
                                       .clkin_from_pll_c0(clkin_from_pll_c0)
                                   );
    defparam           primitive_instance.clkdiv                          = clkdiv;
    defparam           primitive_instance.tsclkdiv                        = tsclkdiv;
    defparam           primitive_instance.tsclksel                        = tsclksel;
    defparam           primitive_instance.prescalar                       = prescalar;
    defparam           primitive_instance.refsel                          = refsel;
    defparam           primitive_instance.device_partname_fivechar_prefix = device_partname_fivechar_prefix;
    defparam           primitive_instance.is_this_first_or_second_adc     = is_this_first_or_second_adc;
    defparam           primitive_instance.analog_input_pin_mask           = analog_input_pin_mask;
    defparam           primitive_instance.pwd                             = hard_pwd;
    defparam           primitive_instance.enable_usr_sim                  = enable_usr_sim;
    defparam           primitive_instance.reference_voltage_sim           = reference_voltage_sim;
    defparam           primitive_instance.simfilename_ch0                 = simfilename_ch0;
    defparam           primitive_instance.simfilename_ch1                 = simfilename_ch1;
    defparam           primitive_instance.simfilename_ch2                 = simfilename_ch2;
    defparam           primitive_instance.simfilename_ch3                 = simfilename_ch3;
    defparam           primitive_instance.simfilename_ch4                 = simfilename_ch4;
    defparam           primitive_instance.simfilename_ch5                 = simfilename_ch5;
    defparam           primitive_instance.simfilename_ch6                 = simfilename_ch6;
    defparam           primitive_instance.simfilename_ch7                 = simfilename_ch7;
    defparam           primitive_instance.simfilename_ch8                 = simfilename_ch8;
    defparam           primitive_instance.simfilename_ch9                 = simfilename_ch9;
    defparam           primitive_instance.simfilename_ch10                = simfilename_ch10;
    defparam           primitive_instance.simfilename_ch11                = simfilename_ch11;
    defparam           primitive_instance.simfilename_ch12                = simfilename_ch12;
    defparam           primitive_instance.simfilename_ch13                = simfilename_ch13;
    defparam           primitive_instance.simfilename_ch14                = simfilename_ch14;
    defparam           primitive_instance.simfilename_ch15                = simfilename_ch15;
    defparam           primitive_instance.simfilename_ch16                = simfilename_ch16;
endmodule

